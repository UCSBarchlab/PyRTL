module toplevel(aes_key, aes_plaintext, aes_ciphertext, clk);
    input[127:0] aes_key;
    input[127:0] aes_plaintext;
    input clk;
    output[127:0] aes_ciphertext;

    wire const2887_0;
    wire[7:0] tmp905;
    wire[31:0] tmp29;
    wire[7:0] tmp1406;
    wire[7:0] tmp240;
    wire[7:0] tmp868;
    wire const1635_0;
    wire[31:0] tmp30;
    wire[7:0] tmp907;
    wire[7:0] tmp241;
    wire[31:0] tmp31;
    wire[255:0] tmp994;
    wire[255:0] tmp2215;
    wire[127:0] temp_25;
    wire[7:0] tmp1639;
    wire[255:0] tmp1633;
    wire[7:0] tmp909;
    wire[255:0] tmp1694;
    wire[247:0] tmp524;
    wire[7:0] tmp242;
    wire[255:0] tmp1055;
    wire[7:0] tmp583;
    wire[7:0] const198_8;
    wire[7:0] tmp910;
    wire[7:0] tmp2396;
    wire const1643_0;
    wire[31:0] tmp33;
    wire[7:0] tmp1795;
    wire[7:0] c1_w39;
    wire[7:0] c2_w39;
    wire[255:0] tmp1642;
    wire[7:0] c3_w39;
    wire[7:0] a1_w7;
    wire[31:0] tmp230;
    wire[247:0] tmp2206;
    wire[7:0] a2_w7;
    wire[7:0] a3_w7;
    wire[255:0] tmp1116;
    wire[127:0] tmp913;
    wire[7:0] tmp34;
    wire[247:0] tmp2467;
    wire[247:0] tmp1644;
    wire[7:0] tmp637;
    wire[127:0] tmp244;
    wire[255:0] tmp1645;
    wire[127:0] tmp892;
    wire[7:0] tmp906;
    wire[31:0] concat_w35;
    wire[7:0] tmp35;
    wire[7:0] tmp915;
    wire[7:0] tmp355;
    wire[255:0] tmp1650;
    wire[127:0] tmp245;
    wire[7:0] tmp2399;
    wire[7:0] tmp916;
    wire[255:0] tmp1384;
    wire[7:0] tmp36;
    wire[247:0] tmp1118;
    wire[255:0] tmp1871;
    wire[7:0] tmp917;
    wire[255:0] tmp1413;
    wire[127:0] tmp246;
    wire[127:0] tmp1182;
    wire[7:0] tmp639;
    wire[7:0] tmp37;
    wire[247:0] tmp1636;
    wire[31:0] tmp247;
    wire[7:0] tmp357;
    wire[255:0] tmp490;
    wire[31:0] shifted_w7;
    wire[7:0] tmp640;
    wire[247:0] tmp2732;
    wire[7:0] tmp920;
    wire[7:0] tmp1728;
    wire[7:0] tmp866;
    wire[31:0] xor_w39;
    wire const2498_0;
    wire[7:0] rc1_w39;
    wire[247:0] tmp2443;
    wire[7:0] tmp921;
    wire[7:0] tmp581;
    wire[7:0] rc3_w39;
    wire[7:0] b2_w7;
    wire[7:0] tmp2402;
    wire[7:0] const248_10;
    wire[255:0] tmp1388;
    wire[7:0] const250_0;
    wire[255:0] tmp1119;
    wire[7:0] tmp39;
    wire[7:0] tmp1507;
    wire[7:0] tmp923;
    wire[255:0] tmp541;
    wire[255:0] tmp2128;
    wire[247:0] tmp998;
    wire[7:0] tmp924;
    wire[7:0] tmp40;
    wire[255:0] tmp1637;
    wire[7:0] const251_0;
    wire[255:0] tmp2533;
    wire const363_0;
    wire[127:0] tmp2352;
    wire[7:0] tmp1699;
    wire[255:0] tmp1284;
    wire[7:0] tmp41;
    wire[7:0] tmp908;
    wire const1868_0;
    wire[127:0] tmp594;
    wire[7:0] tmp1286;
    wire[7:0] tmp927;
    wire[255:0] tmp658;
    wire[7:0] tmp644;
    wire[7:0] tmp42;
    wire[127:0] tmp595;
    wire[255:0] tmp1124;
    wire const1290_0;
    wire[127:0] tmp2354;
    wire[7:0] tmp2382;
    wire[255:0] tmp542;
    wire[7:0] tmp929;
    wire[7:0] c1_w7;
    wire[7:0] tmp645;
    wire[127:0] tmp596;
    wire[7:0] tmp867;
    wire[7:0] tmp930;
    wire[255:0] tmp401;
    wire[7:0] c4_w7;
    wire[7:0] tmp1514;
    wire[7:0] tmp932;
    wire[255:0] tmp1409;
    wire[7:0] tmp933;
    wire[7:0] tmp934;
    wire[7:0] tmp2407;
    wire[7:0] tmp935;
    wire[127:0] tmp2356;
    wire[247:0] tmp1122;
    wire[7:0] tmp937;
    wire[127:0] tmp44;
    wire[7:0] tmp939;
    wire[7:0] tmp940;
    wire[247:0] tmp2760;
    wire[127:0] tmp2357;
    wire[7:0] tmp942;
    wire const375_0;
    wire[31:0] tmp32;
    wire[127:0] tmp45;
    wire[7:0] tmp944;
    wire[247:0] tmp1062;
    wire[7:0] tmp945;
    wire const949_0;
    wire[7:0] tmp648;
    wire[255:0] tmp952;
    wire[127:0] tmp46;
    wire[127:0] tmp600;
    wire const495_0;
    wire[127:0] tmp2068;
    wire[255:0] tmp947;
    wire[247:0] tmp693;
    wire[7:0] tmp649;
    wire[255:0] tmp2216;
    wire[31:0] tmp47;
    wire[127:0] temp_28;
    wire[127:0] tmp601;
    wire[255:0] tmp1305;
    wire[247:0] tmp950;
    wire[31:0] xor_w7;
    wire[7:0] rc1_w7;
    wire const2414_0;
    wire[7:0] rc2_w7;
    wire[247:0] tmp813;
    wire[7:0] rc3_w7;
    wire[7:0] rc4_w7;
    wire[7:0] const48_2;
    wire[255:0] tmp1063;
    wire const953_0;
    wire[247:0] tmp1303;
    wire[255:0] tmp2417;
    wire[255:0] tmp1646;
    wire[255:0] tmp1304;
    wire[31:0] tmp155;
    wire[7:0] tmp605;
    wire[7:0] tmp1511;
    wire[7:0] const51_0;
    wire[7:0] tmp311;
    wire[247:0] tmp1307;
    wire[7:0] tmp911;
    wire[7:0] tmp606;
    wire[7:0] const52_0;
    wire[255:0] tmp2472;
    wire const961_0;
    wire[7:0] tmp607;
    wire[7:0] tmp216;
    wire[255:0] tmp1003;
    wire[31:0] concat_w7;
    wire[255:0] tmp1385;
    wire[31:0] tmp53;
    wire[255:0] tmp498;
    wire[127:0] tmp170;
    wire[7:0] const252_0;
    wire const1422_0;
    wire[7:0] rc3_w27;
    wire[31:0] concat_w39;
    wire[255:0] tmp1007;
    wire const1928_0;
    wire[31:0] tmp253;
    wire[7:0] tmp2091;
    wire[31:0] substituted_w35;
    wire[7:0] tmp2687;
    wire[255:0] tmp2412;
    wire[255:0] tmp2733;
    wire[7:0] tmp1729;
    wire[31:0] tmp254;
    wire[7:0] c4_w39;
    wire[7:0] tmp2688;
    wire const463_0;
    wire[7:0] tmp2689;
    wire[7:0] tmp584;
    wire[7:0] tmp2690;
    wire[127:0] tmp1177;
    wire[31:0] tmp255;
    wire const1832_0;
    wire[255:0] tmp1702;
    wire[7:0] tmp2692;
    wire[31:0] tmp256;
    wire[31:0] substituted_w39;
    wire[7:0] tmp2694;
    wire[31:0] tmp257;
    wire[127:0] tmp1762;
    wire[7:0] tmp2696;
    wire[127:0] tmp554;
    wire[31:0] tmp258;
    wire[247:0] tmp488;
    wire[7:0] tmp2698;
    wire[1407:0] tmp259;
    wire[255:0] tmp372;
    wire[127:0] tmp243;
    wire[7:0] tmp2700;
    wire[7:0] tmp2374;
    wire[7:0] tmp2701;
    wire[127:0] new_2;
    wire[127:0] tmp93;
    wire[7:0] tmp2702;
    wire[7:0] tmp2703;
    wire[255:0] tmp654;
    wire[255:0] tmp778;
    wire[127:0] input_wire_1;
    wire const2217_0;
    wire[255:0] tmp2710;
    wire[7:0] a4_w7;
    wire[255:0] tmp2704;
    wire[127:0] new_1;
    wire[127:0] tmp2648;
    wire[127:0] tmp260;
    wire[255:0] tmp2705;
    wire[247:0] tmp2218;
    wire[127:0] tmp261;
    wire[255:0] tmp1126;
    wire[255:0] tmp2706;
    wire[255:0] tmp1688;
    wire[7:0] tmp2962;
    wire[247:0] tmp2708;
    wire[255:0] tmp2764;
    wire[7:0] tmp262;
    wire[255:0] tmp2283;
    wire[7:0] tmp263;
    wire[7:0] tmp624;
    wire[31:0] tmp188;
    wire const2711_0;
    wire const1009_0;
    wire[247:0] tmp2712;
    wire[31:0] tmp232;
    wire[7:0] tmp264;
    wire[127:0] tmp1472;
    wire[255:0] tmp2713;
    wire[255:0] tmp690;
    wire[7:0] tmp265;
    wire[7:0] tmp137;
    wire[7:0] tmp2715;
    wire[255:0] tmp1268;
    wire[7:0] tmp266;
    wire[127:0] tmp893;
    wire[7:0] tmp914;
    wire[127:0] tmp94;
    wire[7:0] tmp267;
    wire const2719_0;
    wire[247:0] tmp657;
    wire[255:0] tmp2722;
    wire[7:0] tmp268;
    wire[255:0] tmp434;
    wire[7:0] tmp2094;
    wire[7:0] tmp269;
    wire[7:0] tmp2763;
    wire[7:0] tmp608;
    wire[255:0] tmp1419;
    wire[7:0] tmp270;
    wire[255:0] tmp2561;
    wire[247:0] tmp1130;
    wire[31:0] tmp54;
    wire[7:0] tmp271;
    wire[255:0] tmp1317;
    wire[127:0] tmp296;
    wire[7:0] tmp610;
    wire[255:0] tmp1128;
    wire[7:0] tmp272;
    wire const2012_0;
    wire[127:0] tmp2964;
    wire[31:0] tmp56;
    wire[255:0] tmp1240;
    wire[7:0] tmp273;
    wire[255:0] tmp2766;
    wire[31:0] tmp57;
    wire[7:0] c3_w27;
    wire[7:0] tmp612;
    wire[31:0] tmp58;
    wire[247:0] tmp1315;
    wire[127:0] tmp1764;
    wire[7:0] a1_w11;
    wire[7:0] tmp275;
    wire[7:0] a3_w11;
    wire[7:0] a4_w11;
    wire const1647_0;
    wire[7:0] tmp59;
    wire[127:0] temp_16;
    wire[255:0] tmp1321;
    wire[7:0] tmp615;
    wire[7:0] tmp2092;
    wire[7:0] tmp277;
    wire[247:0] tmp2419;
    wire[127:0] input_wire_7;
    wire[247:0] tmp1648;
    wire[7:0] tmp278;
    wire[7:0] tmp279;
    wire const2289_0;
    wire[7:0] tmp141;
    wire[7:0] tmp617;
    wire[255:0] tmp1674;
    wire[255:0] tmp1709;
    wire const1302_0;
    wire[7:0] tmp282;
    wire[127:0] temp_32;
    wire[7:0] tmp2377;
    wire[127:0] tmp2019;
    wire[255:0] tmp1008;
    wire[7:0] tmp285;
    wire[255:0] tmp2802;
    wire[127:0] tmp2378;
    wire[7:0] tmp287;
    wire[255:0] tmp492;
    wire[7:0] tmp1755;
    wire[7:0] tmp288;
    wire[7:0] tmp1730;
    wire[7:0] tmp289;
    wire[247:0] tmp404;
    wire[7:0] tmp2020;
    wire[7:0] tmp291;
    wire[7:0] tmp1236;
    wire[7:0] tmp292;
    wire[7:0] tmp293;
    wire[247:0] tmp661;
    wire const1679_0;
    wire[255:0] tmp1682;
    wire[255:0] tmp1649;
    wire[247:0] tmp1327;
    wire[7:0] b1_w11;
    wire[247:0] tmp2804;
    wire[7:0] b2_w11;
    wire[255:0] tmp1328;
    wire[127:0] tmp295;
    wire[7:0] tmp312;
    wire[7:0] tmp64;
    wire[7:0] tmp2024;
    wire const1330_0;
    wire[7:0] tmp2097;
    wire[247:0] tmp1331;
    wire[7:0] tmp2025;
    wire[7:0] tmp1522;
    wire[7:0] tmp65;
    wire[255:0] tmp1332;
    wire[7:0] tmp2026;
    wire[255:0] tmp1851;
    wire[255:0] tmp493;
    wire[127:0] tmp2651;
    wire[7:0] tmp1334;
    wire const1683_0;
    wire[255:0] tmp662;
    wire[247:0] tmp1684;
    wire[7:0] tmp918;
    wire[7:0] tmp628;
    wire[255:0] tmp1341;
    wire[255:0] tmp2805;
    wire[7:0] const126_0;
    wire[7:0] tmp1234;
    wire[255:0] tmp959;
    wire[7:0] tmp873;
    wire[247:0] tmp1134;
    wire[247:0] tmp2720;
    wire[255:0] tmp960;
    wire[7:0] tmp217;
    wire[127:0] tmp587;
    wire[7:0] tmp571;
    wire[247:0] tmp1708;
    wire[247:0] tmp962;
    wire[7:0] tmp1524;
    wire[7:0] tmp2031;
    wire[127:0] tmp1475;
    wire[255:0] tmp963;
    wire[7:0] tmp2032;
    wire[31:0] tmp113;
    wire[247:0] tmp2724;
    wire[255:0] tmp968;
    wire[255:0] tmp1335;
    wire const965_0;
    wire[255:0] tmp785;
    wire[247:0] tmp966;
    wire[7:0] tmp919;
    wire[7:0] tmp2034;
    wire[31:0] tmp97;
    wire[255:0] tmp967;
    wire[7:0] tmp236;
    wire[7:0] tmp1167;
    wire[7:0] tmp2035;
    wire[7:0] tmp969;
    wire[255:0] tmp1135;
    wire[7:0] tmp2036;
    wire[255:0] tmp827;
    wire[127:0] tmp2652;
    wire[255:0] tmp2734;
    wire[127:0] tmp171;
    wire[7:0] tmp2038;
    wire[255:0] tmp699;
    wire[255:0] tmp2228;
    wire const973_0;
    wire[127:0] temp_34;
    wire[255:0] tmp976;
    wire[255:0] tmp1420;
    wire const1655_0;
    wire[255:0] tmp970;
    wire[247:0] tmp1010;
    wire[7:0] tmp2042;
    wire[7:0] tmp2043;
    wire[255:0] tmp971;
    wire[255:0] tmp2156;
    wire[127:0] tmp299;
    wire[7:0] tmp2045;
    wire[255:0] tmp819;
    wire[7:0] tmp2046;
    wire[255:0] tmp1658;
    wire[255:0] tmp972;
    wire[7:0] tmp1517;
    wire[7:0] tmp2048;
    wire[7:0] tmp2049;
    wire[7:0] tmp2050;
    wire[247:0] tmp2230;
    wire[7:0] tmp2051;
    wire[255:0] tmp975;
    wire[255:0] tmp1652;
    wire[127:0] tmp2052;
    wire[255:0] tmp437;
    wire[247:0] tmp2736;
    wire[255:0] tmp2291;
    wire[255:0] tmp980;
    wire[31:0] tmp158;
    wire const977_0;
    wire[7:0] tmp1171;
    wire[247:0] tmp978;
    wire[255:0] tmp1333;
    wire[127:0] tmp2053;
    wire[127:0] tmp2358;
    wire[247:0] tmp1014;
    wire[255:0] tmp979;
    wire[7:0] rc1_w15;
    wire[7:0] rc1_w27;
    wire[7:0] tmp870;
    wire[7:0] tmp981;
    wire[7:0] rc2_w39;
    wire[255:0] tmp951;
    wire[255:0] tmp2746;
    wire[247:0] tmp1243;
    wire[255:0] tmp2740;
    wire const985_0;
    wire[127:0] tmp1189;
    wire[255:0] tmp988;
    wire[7:0] tmp2799;
    wire[255:0] tmp982;
    wire[255:0] tmp1653;
    wire const2450_0;
    wire[7:0] rc3_w15;
    wire[255:0] tmp983;
    wire[7:0] tmp585;
    wire[247:0] tmp1339;
    wire[247:0] tmp2744;
    wire[7:0] tmp1731;
    wire[255:0] tmp984;
    wire[7:0] rc4_w39;
    wire[255:0] tmp405;
    wire[247:0] tmp805;
    wire const704_0;
    wire[247:0] tmp986;
    wire[255:0] tmp1858;
    wire[7:0] tmp1687;
    wire[7:0] rc4_w27;
    wire[7:0] a3_w39;
    wire[7:0] tmp630;
    wire[7:0] tmp922;
    wire const2747_0;
    wire[247:0] tmp2748;
    wire[7:0] const98_4;
    wire[255:0] tmp992;
    wire const989_0;
    wire[255:0] tmp2236;
    wire[255:0] tmp2749;
    wire[7:0] tmp313;
    wire[7:0] tmp632;
    wire[7:0] b4_w7;
    wire[7:0] tmp2751;
    wire[255:0] tmp701;
    wire[7:0] tmp633;
    wire[31:0] tmp172;
    wire[7:0] const175_0;
    wire[7:0] tmp993;
    wire[7:0] tmp634;
    wire[127:0] tmp249;
    wire[247:0] tmp1692;
    wire[255:0] tmp2758;
    wire[7:0] tmp2103;
    wire[7:0] tmp635;
    wire const997_0;
    wire[127:0] tmp174;
    wire[255:0] tmp1000;
    wire[7:0] tmp636;
    wire[247:0] tmp1656;
    wire[255:0] tmp1698;
    wire[7:0] tmp2961;
    wire const1695_0;
    wire const531_0;
    wire[255:0] tmp1249;
    wire[7:0] const127_0;
    wire[255:0] tmp995;
    wire[7:0] tmp638;
    wire[255:0] tmp823;
    wire[7:0] tmp2400;
    wire[127:0] tmp297;
    wire[255:0] tmp1697;
    wire[7:0] tmp876;
    wire[127:0] input_wire_4;
    wire[7:0] tmp641;
    wire[7:0] tmp2403;
    wire[7:0] tmp2105;
    wire[7:0] tmp643;
    wire[7:0] tmp2405;
    wire[7:0] a4_w39;
    wire[255:0] tmp999;
    wire[7:0] tmp646;
    wire[127:0] tmp1478;
    wire[7:0] tmp647;
    wire[255:0] tmp1004;
    wire[7:0] tmp2106;
    wire[7:0] tmp2410;
    wire[7:0] a1_w27;
    wire[7:0] tmp650;
    wire[127:0] tmp2060;
    wire[7:0] tmp651;
    wire[255:0] tmp786;
    wire[7:0] tmp652;
    wire[255:0] tmp1657;
    wire const656_0;
    wire[31:0] tmp38;
    wire[255:0] tmp659;
    wire[255:0] tmp2812;
    wire[255:0] tmp653;
    wire[255:0] tmp1678;
    wire[7:0] tmp1005;
    wire[255:0] tmp2413;
    wire[127:0] new_4;
    wire[255:0] tmp2770;
    wire[247:0] tmp2415;
    wire[7:0] tmp2108;
    wire[255:0] tmp1705;
    wire[255:0] tmp1012;
    wire[255:0] tmp1357;
    wire[255:0] tmp1006;
    wire[127:0] temp_37;
    wire[255:0] tmp1710;
    wire[31:0] tmp63;
    wire[7:0] tmp325;
    wire const1707_0;
    wire[255:0] tmp1011;
    wire[255:0] tmp2421;
    wire[255:0] tmp534;
    wire[255:0] tmp1248;
    wire const2418_0;
    wire[7:0] tmp856;
    wire[247:0] tmp2768;
    wire[7:0] tmp1238;
    wire[7:0] tmp2237;
    wire[255:0] tmp663;
    wire const660_0;
    wire[7:0] tmp925;
    wire[127:0] tmp1474;
    wire[255:0] tmp2420;
    wire[7:0] tmp1711;
    wire[255:0] tmp1043;
    wire[7:0] const101_0;
    wire[7:0] tmp2422;
    wire[255:0] tmp1272;
    wire const1338_0;
    wire[255:0] tmp1676;
    wire[127:0] tmp2057;
    wire[127:0] tmp1770;
    wire[7:0] a2_w27;
    wire[255:0] tmp1336;
    wire[127:0] tmp2058;
    wire[127:0] tmp1479;
    wire[255:0] tmp1337;
    wire[7:0] a3_w23;
    wire[7:0] tmp2657;
    wire[127:0] tmp300;
    wire[127:0] tmp1185;
    wire[127:0] tmp2059;
    wire[255:0] tmp1340;
    wire[127:0] tmp301;
    wire[255:0] tmp706;
    wire[255:0] tmp1345;
    wire const1342_0;
    wire[7:0] const177_0;
    wire[247:0] tmp1343;
    wire[127:0] temp_38;
    wire[7:0] tmp926;
    wire[127:0] tmp302;
    wire[255:0] tmp1344;
    wire[127:0] tmp2061;
    wire const1242_0;
    wire const2241_0;
    wire[7:0] tmp1346;
    wire[127:0] tmp303;
    wire[7:0] tmp878;
    wire[127:0] tmp2062;
    wire[247:0] tmp2816;
    wire const1350_0;
    wire const1539_0;
    wire[255:0] tmp2481;
    wire[255:0] tmp1353;
    wire[255:0] tmp1347;
    wire[127:0] tmp2063;
    wire[31:0] concat_w15;
    wire[255:0] tmp1348;
    wire[127:0] tmp305;
    wire[31:0] concat_w27;
    wire[31:0] tmp228;
    wire[255:0] tmp1349;
    wire[127:0] tmp1480;
    wire[255:0] tmp1700;
    wire[247:0] tmp1351;
    wire[31:0] xor_w15;
    wire[127:0] tmp306;
    wire[7:0] tmp551;
    wire[255:0] tmp830;
    wire[255:0] tmp1352;
    wire[255:0] tmp2416;
    wire[127:0] tmp307;
    wire[247:0] tmp709;
    wire const1354_0;
    wire[127:0] tmp2066;
    wire[255:0] tmp1361;
    wire[247:0] tmp1423;
    wire[127:0] tmp308;
    wire[127:0] tmp2360;
    wire[127:0] tmp2067;
    wire[7:0] tmp2625;
    wire[7:0] tmp1358;
    wire[127:0] tmp304;
    wire[255:0] tmp818;
    wire[7:0] tmp1732;
    wire[127:0] tmp309;
    wire[7:0] tmp879;
    wire[7:0] tmp928;
    wire[7:0] tmp2381;
    wire[31:0] tmp222;
    wire const1362_0;
    wire[7:0] tmp627;
    wire[255:0] tmp1365;
    wire[255:0] tmp1359;
    wire[255:0] tmp2797;
    wire[247:0] tmp440;
    wire[7:0] tmp2070;
    wire[255:0] tmp710;
    wire[7:0] tmp1157;
    wire[7:0] tmp67;
    wire[7:0] tmp2071;
    wire[255:0] tmp1293;
    wire[255:0] tmp814;
    wire[255:0] tmp1718;
    wire[255:0] tmp1712;
    wire[255:0] tmp1252;
    wire[7:0] c1_w11;
    wire[31:0] xor_w27;
    wire[7:0] c2_w11;
    wire[7:0] tmp1543;
    wire[255:0] tmp1364;
    wire[7:0] c4_w11;
    wire[255:0] tmp1287;
    wire[31:0] substituted_w11;
    wire[247:0] tmp954;
    wire[255:0] tmp1369;
    wire[255:0] tmp1075;
    wire const1366_0;
    wire[247:0] tmp1367;
    wire[255:0] tmp1301;
    wire[7:0] tmp2075;
    wire[127:0] tmp69;
    wire[31:0] xor_w35;
    wire[7:0] tmp317;
    wire[7:0] tmp586;
    wire[7:0] tmp1165;
    wire[255:0] tmp1722;
    wire[31:0] concat_w31;
    wire[127:0] tmp1178;
    wire const1719_0;
    wire[127:0] tmp70;
    wire[7:0] c2_w7;
    wire[255:0] tmp1044;
    wire[7:0] rc1_w35;
    wire[7:0] tmp319;
    wire[255:0] tmp1377;
    wire[31:0] tmp180;
    wire[7:0] tmp1274;
    wire[255:0] tmp1371;
    wire[7:0] tmp1723;
    wire[7:0] c3_w7;
    wire[7:0] tmp2960;
    wire[255:0] tmp1372;
    wire[255:0] tmp2120;
    wire[7:0] tmp1204;
    wire[7:0] tmp321;
    wire[7:0] tmp159;
    wire[31:0] tmp72;
    wire[127:0] tmp2064;
    wire[127:0] tmp1724;
    wire[247:0] tmp1672;
    wire[7:0] tmp322;
    wire[7:0] tmp931;
    wire[255:0] tmp377;
    wire[247:0] tmp1375;
    wire[7:0] b1_w7;
    wire[31:0] xor_w11;
    wire[7:0] rc3_w35;
    wire[7:0] tmp323;
    wire[7:0] tmp604;
    wire[7:0] rc2_w11;
    wire[255:0] tmp833;
    wire[7:0] rc3_w11;
    wire[7:0] tmp324;
    wire[31:0] substituted_w7;
    wire[7:0] const73_3;
    wire[7:0] const75_0;
    wire[7:0] rc4_w35;
    wire[7:0] tmp2084;
    wire[127:0] tmp1726;
    wire[7:0] tmp1818;
    wire[255:0] tmp2223;
    wire[7:0] tmp326;
    wire[127:0] tmp43;
    wire[7:0] rc3_w3;
    wire[7:0] tmp2823;
    wire[127:0] tmp327;
    wire[31:0] tmp204;
    wire[7:0] tmp1166;
    wire[7:0] const76_0;
    wire[31:0] tmp203;
    wire[31:0] tmp182;
    wire[255:0] tmp758;
    wire[127:0] tmp298;
    wire[127:0] tmp597;
    wire[7:0] tmp328;
    wire const471_0;
    wire const1386_0;
    wire[7:0] tmp85;
    wire[7:0] const225_0;
    wire[255:0] tmp1389;
    wire[7:0] tmp329;
    wire[255:0] tmp834;
    wire[31:0] tmp78;
    wire[247:0] tmp1291;
    wire[7:0] tmp330;
    wire[31:0] tmp108;
    wire[7:0] tmp114;
    wire[31:0] tmp79;
    wire[7:0] tmp1159;
    wire[7:0] tmp567;
    wire[7:0] tmp331;
    wire[127:0] tmp2065;
    wire[247:0] tmp1387;
    wire[7:0] tmp1235;
    wire[7:0] tmp936;
    wire[31:0] tmp80;
    wire[255:0] tmp2480;
    wire[247:0] tmp2772;
    wire[31:0] tmp81;
    wire[255:0] tmp1545;
    wire const1013_0;
    wire const2426_0;
    wire[7:0] tmp1484;
    wire[255:0] tmp2754;
    wire[255:0] tmp2429;
    wire[31:0] tmp83;
    wire[7:0] tmp1065;
    wire[255:0] tmp1015;
    wire[7:0] a1_w15;
    wire[7:0] a1_w31;
    wire[255:0] tmp2424;
    wire[7:0] a3_w15;
    wire[7:0] tmp938;
    wire[7:0] a4_w15;
    wire[255:0] tmp2425;
    wire const1414_0;
    wire[255:0] tmp2782;
    wire[7:0] tmp629;
    wire[247:0] tmp2427;
    wire[7:0] a2_w31;
    wire const1021_0;
    wire[255:0] tmp1024;
    wire[127:0] tmp598;
    wire[255:0] tmp1018;
    wire[255:0] tmp474;
    wire[7:0] tmp1738;
    wire[255:0] tmp2473;
    wire[255:0] tmp1019;
    wire[7:0] a3_w31;
    wire[7:0] tmp235;
    wire[7:0] tmp1739;
    wire[7:0] tmp86;
    wire[255:0] tmp1020;
    wire[255:0] tmp441;
    wire[7:0] tmp1740;
    wire[7:0] a3_w19;
    wire[247:0] tmp1022;
    wire[247:0] tmp1355;
    wire[7:0] tmp87;
    wire[7:0] tmp2434;
    wire[7:0] tmp941;
    wire const2783_0;
    wire[7:0] b3_w7;
    wire[7:0] a4_w23;
    wire[7:0] tmp1742;
    wire[247:0] tmp2475;
    wire[7:0] tmp556;
    wire[255:0] tmp1028;
    wire[31:0] shifted_w15;
    wire[7:0] tmp184;
    wire[31:0] tmp88;
    wire const2755_0;
    wire[7:0] tmp1744;
    wire const1294_0;
    wire[7:0] tmp1745;
    wire[255:0] tmp1027;
    wire[255:0] tmp370;
    wire[7:0] b1_w15;
    wire[7:0] b2_w15;
    wire[255:0] tmp838;
    wire[7:0] b3_w15;
    wire[7:0] b4_w15;
    wire[7:0] tmp943;
    wire const2791_0;
    wire[255:0] tmp469;
    wire[255:0] tmp2794;
    wire[255:0] tmp1072;
    wire[7:0] tmp1753;
    wire[7:0] tmp161;
    wire const1033_0;
    wire[255:0] tmp1356;
    wire[255:0] tmp1036;
    wire[7:0] tmp1756;
    wire[127:0] tmp599;
    wire[7:0] tmp1757;
    wire[255:0] tmp1906;
    wire[7:0] tmp1758;
    wire[247:0] tmp368;
    wire[255:0] tmp1031;
    wire const2442_0;
    wire[7:0] tmp190;
    wire[247:0] tmp2792;
    wire[255:0] tmp1032;
    wire[255:0] tmp2793;
    wire[247:0] tmp1584;
    wire[127:0] tmp1760;
    wire[7:0] tmp92;
    wire[7:0] tmp2446;
    wire const2795_0;
    wire const2538_0;
    wire[247:0] tmp2439;
    wire[247:0] tmp2796;
    wire[255:0] tmp1040;
    wire[7:0] c1_w15;
    wire[7:0] c2_w15;
    wire[7:0] tmp2096;
    wire const840_0;
    wire[127:0] tmp218;
    wire[7:0] tmp2044;
    wire[7:0] tmp844;
    wire[255:0] tmp1838;
    wire[255:0] tmp1874;
    wire[7:0] tmp664;
    wire[255:0] tmp369;
    wire[127:0] tmp2055;
    wire const2253_0;
    wire[7:0] tmp2225;
    wire const824_0;
    wire[255:0] tmp946;
    wire const668_0;
    wire[255:0] tmp1300;
    wire[255:0] tmp671;
    wire[255:0] tmp1585;
    wire[255:0] tmp665;
    wire[127:0] tmp891;
    wire[7:0] tmp1169;
    wire[255:0] tmp2256;
    wire[255:0] tmp666;
    wire[7:0] tmp1298;
    wire[255:0] tmp2509;
    wire[255:0] tmp667;
    wire[247:0] tmp1552;
    wire[247:0] tmp669;
    wire[255:0] tmp1395;
    wire[255:0] tmp1839;
    wire const1844_0;
    wire[255:0] tmp670;
    wire[7:0] tmp371;
    wire[255:0] tmp675;
    wire[255:0] tmp790;
    wire const672_0;
    wire[127:0] tmp2359;
    wire[247:0] tmp673;
    wire[255:0] tmp1590;
    wire[255:0] tmp674;
    wire[7:0] tmp1489;
    wire[7:0] tmp676;
    wire[247:0] tmp1070;
    wire[255:0] tmp1553;
    wire const680_0;
    wire[7:0] tmp341;
    wire[255:0] tmp683;
    wire[255:0] tmp1689;
    wire[255:0] tmp677;
    wire[247:0] tmp1588;
    wire[7:0] tmp1137;
    wire[7:0] tmp1170;
    wire[7:0] tmp2069;
    wire[255:0] tmp678;
    wire[7:0] tmp1734;
    wire[255:0] tmp948;
    wire[255:0] tmp679;
    wire[247:0] tmp681;
    wire[127:0] tmp1481;
    wire[7:0] tmp1490;
    wire[255:0] tmp682;
    wire[7:0] tmp443;
    wire[255:0] tmp1071;
    wire const1611_0;
    wire[255:0] tmp687;
    wire[7:0] tmp1555;
    wire const684_0;
    wire[255:0] tmp1273;
    wire[247:0] tmp685;
    wire[255:0] tmp1299;
    wire[255:0] tmp1589;
    wire[7:0] tmp557;
    wire[255:0] tmp686;
    wire[255:0] tmp1360;
    wire[7:0] tmp688;
    wire[247:0] tmp532;
    wire[255:0] tmp2131;
    wire[31:0] substituted_w23;
    wire[7:0] tmp332;
    wire[255:0] tmp2447;
    wire[255:0] tmp1039;
    wire[7:0] tmp1491;
    wire[7:0] tmp333;
    wire[255:0] tmp2448;
    wire[255:0] tmp1076;
    wire[7:0] tmp1041;
    wire const1390_0;
    wire[255:0] tmp1878;
    wire[255:0] tmp2449;
    wire[127:0] tmp602;
    wire[247:0] tmp2451;
    wire const1045_0;
    wire[7:0] tmp1591;
    wire[255:0] tmp1048;
    wire[7:0] tmp336;
    wire[255:0] tmp494;
    wire[7:0] tmp1394;
    wire[127:0] tmp168;
    wire[247:0] tmp793;
    wire[31:0] tmp156;
    wire[255:0] tmp2457;
    wire const2454_0;
    wire[255:0] tmp373;
    wire[7:0] tmp115;
    wire const1398_0;
    wire const1715_0;
    wire[255:0] tmp1401;
    wire[247:0] tmp1046;
    wire[7:0] tmp339;
    wire[255:0] tmp1047;
    wire[7:0] tmp2370;
    wire[7:0] tmp340;
    wire[7:0] tmp2929;
    wire[255:0] tmp1052;
    wire[255:0] tmp956;
    wire const1049_0;
    wire[255:0] tmp1875;
    wire[247:0] tmp1050;
    wire[31:0] shifted_w19;
    wire[255:0] tmp2465;
    wire[255:0] tmp2459;
    wire[247:0] tmp1363;
    wire[255:0] tmp1051;
    wire[7:0] const50_0;
    wire[7:0] tmp343;
    wire[7:0] tmp1053;
    wire[255:0] tmp374;
    wire const1402_0;
    wire[7:0] tmp344;
    wire[7:0] tmp2072;
    wire[7:0] tmp345;
    wire[7:0] tmp346;
    wire[127:0] tmp49;
    wire[7:0] tmp347;
    wire[255:0] tmp987;
    wire[255:0] tmp1060;
    wire[255:0] tmp1942;
    wire[255:0] tmp1054;
    wire[7:0] tmp350;
    wire[255:0] tmp497;
    wire[7:0] tmp351;
    wire[7:0] tmp352;
    wire[255:0] tmp1396;
    wire[7:0] tmp353;
    wire[7:0] tmp354;
    wire[247:0] tmp376;
    wire[255:0] tmp1056;
    wire[7:0] tmp356;
    wire[7:0] c3_w11;
    wire[247:0] tmp1058;
    wire[7:0] tmp358;
    wire[255:0] tmp2545;
    wire[7:0] tmp359;
    wire[255:0] tmp1059;
    wire[255:0] tmp1429;
    wire[255:0] tmp366;
    wire[255:0] tmp360;
    wire[7:0] tmp314;
    wire[255:0] tmp1064;
    wire const1061_0;
    wire[255:0] tmp955;
    wire[255:0] tmp361;
    wire[255:0] tmp2477;
    wire const1426_0;
    wire[255:0] tmp2471;
    wire[7:0] a4_w35;
    wire[255:0] tmp362;
    wire[255:0] tmp1309;
    wire[247:0] tmp364;
    wire[7:0] a3_w27;
    wire[7:0] c3_w15;
    wire[7:0] b2_w19;
    wire[7:0] c4_w15;
    wire[7:0] tmp162;
    wire const692_0;
    wire[127:0] tmp68;
    wire[255:0] tmp695;
    wire[255:0] tmp689;
    wire[31:0] tmp13;
    wire[7:0] tmp2093;
    wire const2137_0;
    wire[127:0] tmp1763;
    wire[255:0] tmp2806;
    wire[7:0] tmp574;
    wire[7:0] tmp315;
    wire[255:0] tmp2800;
    wire[255:0] tmp691;
    wire[7:0] tmp957;
    wire[255:0] tmp1846;
    wire const1880_0;
    wire[255:0] tmp2801;
    wire[247:0] tmp2138;
    wire[127:0] tmp95;
    wire[247:0] tmp1716;
    wire[255:0] tmp694;
    wire[255:0] tmp747;
    wire const1306_0;
    wire[127:0] tmp1765;
    wire[127:0] tmp96;
    wire[7:0] tmp503;
    wire[255:0] tmp382;
    wire const696_0;
    wire[247:0] tmp697;
    wire[127:0] tmp219;
    wire[7:0] tmp2098;
    wire[127:0] tmp1766;
    wire[255:0] tmp698;
    wire[247:0] tmp1877;
    wire[7:0] tmp2099;
    wire const379_0;
    wire[247:0] tmp2808;
    wire[127:0] tmp2056;
    wire[7:0] tmp700;
    wire[7:0] tmp316;
    wire[7:0] tmp2100;
    wire const2229_0;
    wire[255:0] tmp2809;
    wire[7:0] tmp2365;
    wire[7:0] rc2_w15;
    wire[7:0] tmp2101;
    wire[127:0] input_wire_11;
    wire[255:0] tmp1078;
    wire[7:0] rc4_w15;
    wire[7:0] tmp274;
    wire[255:0] tmp707;
    wire[255:0] tmp1368;
    wire[7:0] const100_0;
    wire const764_0;
    wire[127:0] tmp99;
    wire[7:0] tmp1784;
    wire[7:0] tmp2104;
    wire[255:0] tmp702;
    wire[247:0] tmp1596;
    wire[127:0] tmp1769;
    wire[7:0] tmp2107;
    wire const1888_0;
    wire[255:0] tmp703;
    wire[7:0] tmp2109;
    wire[255:0] tmp1308;
    wire[255:0] tmp2813;
    wire[247:0] tmp1881;
    wire[7:0] tmp2111;
    wire[7:0] tmp2112;
    wire[7:0] tmp2113;
    wire[7:0] tmp2076;
    wire[7:0] tmp2114;
    wire[255:0] tmp2773;
    wire[7:0] tmp2115;
    wire[255:0] tmp964;
    wire[255:0] tmp711;
    wire const708_0;
    wire[255:0] tmp1079;
    wire const2121_0;
    wire[255:0] tmp2124;
    wire[7:0] tmp1370;
    wire[255:0] tmp2118;
    wire[31:0] tmp104;
    wire[255:0] tmp958;
    wire const2819_0;
    wire[255:0] tmp2119;
    wire[255:0] tmp1597;
    wire[7:0] tmp712;
    wire[31:0] tmp105;
    wire[127:0] tmp1773;
    wire[255:0] tmp2232;
    wire[31:0] tmp106;
    wire[7:0] tmp1310;
    wire[255:0] tmp1428;
    wire[247:0] tmp2122;
    wire const716_0;
    wire[255:0] tmp719;
    wire[127:0] tmp1138;
    wire[255:0] tmp713;
    wire[7:0] tmp318;
    wire[255:0] tmp2741;
    wire[7:0] tmp61;
    wire[255:0] tmp1417;
    wire[7:0] a1_w19;
    wire[7:0] tmp625;
    wire[7:0] a2_w19;
    wire[7:0] tmp383;
    wire const2125_0;
    wire[247:0] tmp2126;
    wire[255:0] tmp1886;
    wire[7:0] tmp109;
    wire const367_0;
    wire[255:0] tmp417;
    wire[255:0] tmp2127;
    wire[7:0] tmp1418;
    wire[255:0] tmp1602;
    wire[255:0] tmp2204;
    wire[127:0] tmp2604;
    wire[7:0] tmp110;
    wire const2478_0;
    wire[247:0] tmp2479;
    wire[7:0] tmp849;
    wire[255:0] tmp1068;
    wire[255:0] tmp1425;
    wire[247:0] tmp1082;
    wire const2133_0;
    wire[255:0] tmp2136;
    wire const1374_0;
    wire[255:0] tmp2130;
    wire[7:0] tmp2482;
    wire[7:0] tmp2685;
    wire[255:0] tmp378;
    wire[7:0] tmp112;
    wire[247:0] tmp1600;
    wire[255:0] tmp1421;
    wire[7:0] tmp280;
    wire const1073_0;
    wire[255:0] tmp504;
    wire[247:0] tmp1074;
    wire[255:0] tmp2489;
    wire[7:0] tmp419;
    wire[247:0] tmp2134;
    wire[7:0] tmp1190;
    wire[255:0] tmp1424;
    wire[127:0] input_wire_5;
    wire[255:0] tmp2737;
    wire[255:0] tmp2135;
    wire[127:0] tmp71;
    wire[255:0] tmp1244;
    wire[7:0] tmp1077;
    wire[7:0] b1_w19;
    wire[127:0] tmp882;
    wire[247:0] tmp1427;
    wire[7:0] tmp2385;
    wire[7:0] b3_w19;
    wire const387_0;
    wire[7:0] b4_w19;
    wire const1081_0;
    wire[7:0] tmp320;
    wire[255:0] tmp1084;
    wire[247:0] tmp380;
    wire[247:0] tmp769;
    wire[7:0] tmp1430;
    wire[255:0] tmp1601;
    wire[255:0] tmp381;
    wire const2490_0;
    wire[247:0] tmp2491;
    wire[255:0] tmp1080;
    wire[7:0] tmp898;
    wire[7:0] tmp116;
    wire[255:0] tmp384;
    wire[255:0] tmp2148;
    wire[255:0] tmp2142;
    wire[255:0] tmp1083;
    wire[255:0] tmp390;
    wire[255:0] tmp2288;
    wire[7:0] tmp117;
    wire[255:0] tmp1088;
    wire[127:0] tmp1432;
    wire const1085_0;
    wire[255:0] tmp385;
    wire[7:0] tmp2080;
    wire[127:0] tmp1433;
    wire[255:0] tmp2774;
    wire[247:0] tmp2146;
    wire[255:0] tmp770;
    wire[7:0] c2_w19;
    wire[7:0] tmp1496;
    wire[7:0] c3_w19;
    wire[7:0] tmp1603;
    wire[7:0] c4_w19;
    wire[7:0] tmp2027;
    wire[7:0] tmp857;
    wire[31:0] substituted_w19;
    wire[127:0] tmp118;
    wire[255:0] tmp389;
    wire[255:0] tmp426;
    wire const2149_0;
    wire[7:0] tmp1435;
    wire[247:0] tmp1086;
    wire[255:0] tmp2274;
    wire[255:0] tmp1373;
    wire[7:0] tmp237;
    wire[255:0] tmp714;
    wire[247:0] tmp2880;
    wire[255:0] tmp2830;
    wire[255:0] tmp2824;
    wire[255:0] tmp2501;
    wire[255:0] tmp715;
    wire[255:0] tmp2476;
    wire[247:0] tmp508;
    wire[255:0] tmp2825;
    wire[255:0] tmp1573;
    wire[7:0] tmp2362;
    wire[255:0] tmp718;
    wire[7:0] c1_w19;
    wire[247:0] tmp2828;
    wire const1892_0;
    wire[255:0] tmp723;
    wire const720_0;
    wire[247:0] tmp721;
    wire[255:0] tmp809;
    wire[7:0] tmp1779;
    wire[255:0] tmp386;
    wire[255:0] tmp722;
    wire[7:0] tmp1780;
    wire[247:0] tmp2832;
    wire[255:0] tmp2180;
    wire[7:0] tmp724;
    wire[7:0] tmp1781;
    wire[127:0] tmp2965;
    wire[255:0] tmp1954;
    wire[255:0] tmp2833;
    wire[7:0] rc1_w11;
    wire[31:0] tmp207;
    wire[7:0] tmp1782;
    wire const728_0;
    wire[7:0] tmp2691;
    wire[255:0] tmp731;
    wire[255:0] tmp725;
    wire[247:0] tmp388;
    wire[127:0] tmp591;
    wire[255:0] tmp1376;
    wire[255:0] tmp726;
    wire[255:0] tmp2842;
    wire[255:0] tmp2836;
    wire[255:0] tmp727;
    wire[7:0] tmp1089;
    wire[247:0] tmp729;
    wire[255:0] tmp2728;
    wire[7:0] tmp1786;
    wire[127:0] tmp590;
    wire const776_0;
    wire[255:0] tmp730;
    wire[7:0] tmp1813;
    wire[7:0] tmp1787;
    wire[7:0] tmp1434;
    wire[247:0] tmp2840;
    wire[255:0] tmp735;
    wire[7:0] tmp2083;
    wire const1057_0;
    wire const732_0;
    wire[247:0] tmp733;
    wire[7:0] tmp1789;
    wire[255:0] tmp2152;
    wire[255:0] tmp734;
    wire const2843_0;
    wire[255:0] tmp1381;
    wire[7:0] tmp1790;
    wire[7:0] tmp736;
    wire[247:0] tmp825;
    wire[247:0] tmp424;
    wire[7:0] tmp1791;
    wire[7:0] tmp2578;
    wire const1378_0;
    wire const740_0;
    wire[255:0] tmp743;
    wire[255:0] tmp737;
    wire[7:0] tmp2386;
    wire[247:0] tmp2150;
    wire[7:0] const201_0;
    wire[7:0] tmp1793;
    wire[255:0] tmp1654;
    wire[255:0] tmp738;
    wire[247:0] tmp1379;
    wire[255:0] tmp2854;
    wire[7:0] tmp1794;
    wire[7:0] tmp2697;
    wire const2546_0;
    wire[255:0] tmp394;
    wire[127:0] tmp119;
    wire[247:0] tmp392;
    wire[255:0] tmp425;
    wire[255:0] tmp393;
    wire[7:0] tmp1453;
    wire[127:0] tmp120;
    wire[255:0] tmp2484;
    wire[247:0] tmp2503;
    wire[7:0] tmp395;
    wire const2157_0;
    wire[7:0] tmp2699;
    wire[7:0] tmp1439;
    wire[255:0] tmp2154;
    wire[1407:0] expanded_key;
    wire[7:0] tmp2506;
    wire[255:0] tmp402;
    wire[255:0] tmp1380;
    wire[255:0] tmp2155;
    wire[31:0] tmp122;
    wire[247:0] tmp2186;
    wire[7:0] tmp1441;
    wire[7:0] tmp1497;
    wire[255:0] tmp397;
    wire const2827_0;
    wire[255:0] tmp2513;
    wire[255:0] tmp1042;
    wire[247:0] tmp2158;
    wire[7:0] rc1_w19;
    wire[7:0] rc2_w19;
    wire[255:0] tmp430;
    wire[7:0] tmp1443;
    wire[7:0] rc4_w19;
    wire[31:0] w1;
    wire[7:0] const123_5;
    wire[7:0] tmp1444;
    wire[255:0] tmp1903;
    wire[127:0] tmp124;
    wire[7:0] a2_w39;
    wire[247:0] tmp2511;
    wire[255:0] tmp406;
    wire[247:0] tmp829;
    wire const403_0;
    wire[31:0] w2;
    wire[7:0] tmp1205;
    wire[255:0] tmp2512;
    wire[7:0] tmp1446;
    wire[7:0] tmp1382;
    wire[255:0] tmp2140;
    wire[7:0] tmp2165;
    wire[255:0] tmp2885;
    wire const2514_0;
    wire[7:0] tmp2363;
    wire[247:0] tmp2515;
    wire[7:0] const102_0;
    wire[7:0] tmp1448;
    wire[7:0] tmp2086;
    wire const2169_0;
    wire[255:0] tmp2172;
    wire const2707_0;
    wire[7:0] tmp1449;
    wire[255:0] tmp1392;
    wire const411_0;
    wire[7:0] const226_0;
    wire[255:0] tmp414;
    wire[255:0] tmp1628;
    wire[255:0] tmp2167;
    wire[31:0] tmp129;
    wire[7:0] tmp1452;
    wire[255:0] tmp2810;
    wire[255:0] tmp409;
    wire[7:0] tmp1454;
    wire[247:0] tmp717;
    wire[31:0] tmp130;
    wire[7:0] tmp631;
    wire[255:0] tmp410;
    wire[247:0] tmp1247;
    wire[31:0] tmp131;
    wire[247:0] tmp412;
    wire[7:0] tmp2189;
    wire[31:0] tmp132;
    wire[7:0] tmp1460;
    wire[7:0] tmp455;
    wire[255:0] tmp413;
    wire[7:0] tmp1462;
    wire[7:0] tmp2087;
    wire[7:0] tmp1212;
    wire[7:0] a1_w23;
    wire[255:0] tmp418;
    wire const415_0;
    wire const1852_0;
    wire[247:0] tmp416;
    wire[7:0] const227_0;
    wire[7:0] tmp134;
    wire[7:0] tmp2074;
    wire const1093_0;
    wire[7:0] tmp851;
    wire[7:0] tmp2634;
    wire[255:0] tmp1096;
    wire[7:0] tmp1455;
    wire[247:0] tmp741;
    wire[7:0] tmp1777;
    wire[7:0] tmp135;
    wire[255:0] tmp516;
    wire[255:0] tmp1091;
    wire[7:0] tmp1735;
    wire[7:0] tmp2129;
    wire[7:0] tmp431;
    wire[7:0] tmp136;
    wire[31:0] tmp6;
    wire const744_0;
    wire[247:0] tmp1660;
    wire[247:0] tmp1094;
    wire[7:0] tmp2088;
    wire[247:0] tmp705;
    wire[247:0] tmp496;
    wire[255:0] tmp826;
    wire const2807_0;
    wire[255:0] tmp746;
    wire[7:0] tmp2388;
    wire[127:0] tmp2932;
    wire[7:0] a2_w23;
    wire[255:0] tmp1100;
    wire const1097_0;
    wire[247:0] tmp1098;
    wire const2193_0;
    wire[31:0] tmp138;
    wire[7:0] tmp2387;
    wire[255:0] tmp2826;
    wire[7:0] tmp1778;
    wire[255:0] tmp1099;
    wire[255:0] tmp755;
    wire[255:0] tmp517;
    wire[255:0] tmp749;
    wire[31:0] shifted_w39;
    wire[7:0] tmp1101;
    wire[7:0] b3_w23;
    wire[255:0] tmp750;
    wire[255:0] tmp2444;
    wire[7:0] tmp139;
    wire[7:0] tmp2089;
    wire[255:0] tmp751;
    wire const2779_0;
    wire[247:0] tmp753;
    wire[7:0] tmp140;
    wire[255:0] tmp1067;
    wire[255:0] tmp2829;
    wire[255:0] tmp2485;
    wire[255:0] tmp754;
    wire const1314_0;
    wire[255:0] tmp782;
    wire[255:0] tmp1104;
    wire const756_0;
    wire[31:0] tmp8;
    wire[247:0] tmp1106;
    wire[7:0] tmp142;
    wire[255:0] tmp438;
    wire[127:0] tmp1431;
    wire[255:0] tmp1967;
    wire[255:0] tmp1112;
    wire[127:0] tmp1139;
    wire[7:0] tmp1250;
    wire const1109_0;
    wire[7:0] b1_w27;
    wire[7:0] tmp2090;
    wire[7:0] a2_w35;
    wire[247:0] tmp1110;
    wire[7:0] c2_w23;
    wire[255:0] tmp432;
    wire[7:0] c3_w23;
    wire[7:0] c4_w23;
    wire[255:0] tmp2834;
    wire[255:0] tmp797;
    wire[255:0] tmp767;
    wire[127:0] tmp592;
    wire[255:0] tmp761;
    wire[255:0] tmp1907;
    wire[7:0] c1_w31;
    wire[7:0] tmp1113;
    wire[31:0] tmp238;
    wire[255:0] tmp1280;
    wire[255:0] tmp1717;
    wire[255:0] tmp2709;
    wire[255:0] tmp762;
    wire const2831_0;
    wire const1948_0;
    wire[127:0] tmp144;
    wire[255:0] tmp763;
    wire[255:0] tmp1120;
    wire[247:0] tmp765;
    wire[127:0] tmp1768;
    wire[7:0] tmp2364;
    wire[127:0] tmp145;
    wire[255:0] tmp1023;
    wire[255:0] tmp1115;
    wire[127:0] tmp221;
    wire[255:0] tmp2849;
    wire[255:0] tmp1264;
    wire[255:0] tmp2192;
    wire[127:0] tmp1467;
    wire[127:0] tmp2085;
    wire[7:0] tmp1796;
    wire const2771_0;
    wire[247:0] tmp2852;
    wire[127:0] tmp1468;
    wire[255:0] tmp2714;
    wire[7:0] tmp349;
    wire[31:0] tmp28;
    wire[255:0] tmp2853;
    wire[7:0] a2_w3;
    wire[7:0] tmp1798;
    wire const2185_0;
    wire[7:0] tmp2029;
    wire const1121_0;
    wire[127:0] tmp845;
    wire[127:0] tmp1469;
    wire const1988_0;
    wire const2855_0;
    wire[247:0] tmp2856;
    wire[255:0] tmp1123;
    wire[7:0] tmp611;
    wire[31:0] tmp231;
    wire[7:0] tmp1800;
    wire[255:0] tmp2857;
    wire[255:0] tmp1016;
    wire[7:0] tmp1125;
    wire[7:0] tmp1801;
    wire const788_0;
    wire[7:0] tmp2859;
    wire[7:0] tmp1502;
    wire[7:0] tmp1802;
    wire const1129_0;
    wire[7:0] tmp1733;
    wire[255:0] tmp1132;
    wire[7:0] tmp1803;
    wire[7:0] tmp852;
    wire[255:0] tmp2866;
    wire[7:0] tmp1458;
    wire[255:0] tmp2860;
    wire[7:0] tmp9;
    wire[247:0] tmp2487;
    wire[7:0] tmp1804;
    wire[31:0] tmp103;
    wire[255:0] tmp2568;
    wire[31:0] tmp82;
    wire[255:0] tmp2861;
    wire[7:0] tmp1805;
    wire[247:0] tmp436;
    wire[127:0] tmp1473;
    wire[31:0] w5;
    wire[255:0] tmp2862;
    wire[7:0] tmp2835;
    wire[7:0] tmp1806;
    wire[247:0] tmp2864;
    wire[127:0] input_wire_3;
    wire[255:0] tmp1131;
    wire[7:0] tmp1807;
    wire[255:0] tmp2865;
    wire[255:0] tmp1136;
    wire[127:0] tmp894;
    wire[7:0] tmp1808;
    wire[255:0] tmp2870;
    wire[255:0] tmp2423;
    wire const2867_0;
    wire[247:0] tmp2868;
    wire[7:0] tmp1810;
    wire[7:0] tmp1811;
    wire[7:0] tmp1783;
    wire[255:0] tmp2869;
    wire[127:0] tmp1476;
    wire const2305_0;
    wire[7:0] tmp2775;
    wire[7:0] c3_w31;
    wire[7:0] tmp1814;
    wire[7:0] tmp1815;
    wire[127:0] tmp2896;
    wire[247:0] tmp1403;
    wire[7:0] tmp1816;
    wire[7:0] tmp1817;
    wire[255:0] tmp420;
    wire[7:0] a1_w39;
    wire[127:0] tmp1477;
    wire[7:0] tmp1819;
    wire[127:0] new_3;
    wire[255:0] tmp2139;
    wire[7:0] tmp1820;
    wire[255:0] tmp2716;
    wire[7:0] tmp1821;
    wire[7:0] tmp1822;
    wire[7:0] tmp901;
    wire[7:0] tmp1823;
    wire const1972_0;
    wire[7:0] tmp1824;
    wire[255:0] tmp1634;
    wire const1828_0;
    wire[7:0] a2_w15;
    wire[255:0] tmp1831;
    wire[255:0] tmp1825;
    wire[255:0] tmp533;
    wire[255:0] tmp2529;
    wire const2839_0;
    wire const2526_0;
    wire[255:0] tmp1826;
    wire[7:0] tmp1017;
    wire[127:0] tmp146;
    wire[255:0] tmp442;
    wire[255:0] tmp1827;
    wire[7:0] tmp2315;
    wire[247:0] tmp1829;
    wire[7:0] tmp2530;
    wire[7:0] b4_w27;
    wire const1912_0;
    wire[31:0] tmp147;
    wire[255:0] tmp1830;
    wire const439_0;
    wire[7:0] a2_w11;
    wire const2534_0;
    wire[255:0] tmp1312;
    wire[255:0] tmp1114;
    wire[255:0] tmp2537;
    wire[7:0] tmp84;
    wire[7:0] rc2_w23;
    wire[255:0] tmp1285;
    wire[7:0] rc3_w23;
    wire[247:0] tmp789;
    wire[7:0] rc4_w23;
    wire[7:0] const148_6;
    wire[7:0] tmp1785;
    wire[7:0] const150_0;
    wire[127:0] tmp149;
    wire[255:0] tmp1909;
    wire[7:0] tmp1836;
    wire[247:0] tmp2535;
    wire[7:0] tmp1485;
    wire[255:0] tmp1970;
    wire[7:0] tmp2371;
    wire[255:0] tmp2536;
    wire[255:0] tmp2776;
    wire[7:0] tmp2102;
    wire[255:0] tmp1843;
    wire[255:0] tmp1837;
    wire[255:0] tmp2541;
    wire[7:0] tmp1487;
    wire[255:0] tmp2837;
    wire[247:0] tmp2539;
    wire[7:0] tmp1737;
    wire[7:0] tmp1488;
    wire[255:0] tmp2540;
    wire[7:0] tmp2201;
    wire[7:0] tmp2871;
    wire[247:0] tmp1841;
    wire[7:0] tmp479;
    wire[255:0] tmp2440;
    wire[7:0] tmp2542;
    wire[31:0] tmp154;
    wire[127:0] tmp1187;
    wire[255:0] tmp1842;
    wire[255:0] tmp2750;
    wire[7:0] tmp1486;
    wire[255:0] tmp1847;
    wire[7:0] tmp897;
    wire[255:0] tmp1971;
    wire[255:0] tmp2549;
    wire[255:0] tmp1662;
    wire[247:0] tmp1845;
    wire[255:0] tmp2428;
    wire[31:0] substituted_w31;
    wire[7:0] tmp1492;
    wire[31:0] tmp157;
    wire[255:0] tmp2544;
    wire[7:0] tmp1493;
    wire[7:0] tmp1503;
    wire[255:0] tmp2838;
    wire[255:0] tmp1030;
    wire[7:0] tmp1848;
    wire[7:0] tmp2607;
    wire[127:0] tmp2946;
    wire[7:0] tmp1494;
    wire[247:0] tmp2547;
    wire[255:0] tmp2777;
    wire[255:0] tmp2717;
    wire[7:0] a4_w27;
    wire[7:0] tmp1495;
    wire[7:0] tmp12;
    wire[255:0] tmp2488;
    wire[255:0] tmp2548;
    wire[7:0] tmp1223;
    wire[255:0] tmp1855;
    wire[255:0] tmp1849;
    wire[127:0] tmp2018;
    wire[255:0] tmp2553;
    wire[7:0] tmp160;
    wire[255:0] tmp1850;
    wire[127:0] tmp1499;
    wire[255:0] tmp2433;
    wire[31:0] xor_w3;
    wire[255:0] tmp766;
    wire[247:0] tmp2876;
    wire[255:0] tmp771;
    wire const768_0;
    wire[127:0] tmp1188;
    wire const2181_0;
    wire[255:0] tmp2184;
    wire const1659_0;
    wire[255:0] tmp2178;
    wire const423_0;
    wire[7:0] tmp1788;
    wire const2879_0;
    wire[127:0] tmp593;
    wire[255:0] tmp2179;
    wire[247:0] tmp2431;
    wire[127:0] tmp193;
    wire[7:0] tmp772;
    wire[7:0] b2_w39;
    wire[247:0] tmp1720;
    wire[247:0] tmp2009;
    wire[255:0] tmp2881;
    wire[255:0] tmp2841;
    wire[247:0] tmp2182;
    wire[7:0] tmp2883;
    wire[255:0] tmp1641;
    wire[255:0] tmp779;
    wire[255:0] tmp773;
    wire[247:0] tmp1026;
    wire[255:0] tmp2188;
    wire[7:0] tmp563;
    wire[255:0] tmp2890;
    wire[7:0] tmp850;
    wire[7:0] tmp1191;
    wire[255:0] tmp2884;
    wire[255:0] tmp775;
    wire[7:0] tmp609;
    wire[255:0] tmp2468;
    wire const427_0;
    wire[255:0] tmp2187;
    wire[255:0] tmp1979;
    wire[255:0] tmp2781;
    wire[255:0] tmp2886;
    wire[7:0] tmp1809;
    wire[247:0] tmp1889;
    wire[255:0] tmp1661;
    wire[7:0] tmp2811;
    wire[247:0] tmp2888;
    wire[255:0] tmp783;
    wire[255:0] tmp2846;
    wire const780_0;
    wire[255:0] tmp2889;
    wire[255:0] tmp2196;
    wire[255:0] tmp2190;
    wire[255:0] tmp444;
    wire[255:0] tmp2894;
    wire const2891_0;
    wire[247:0] tmp1977;
    wire[255:0] tmp2191;
    wire[7:0] tmp784;
    wire[7:0] tmp1741;
    wire[7:0] b3_w39;
    wire[255:0] tmp2893;
    wire[255:0] tmp1311;
    wire[255:0] tmp2543;
    wire[7:0] tmp2367;
    wire[247:0] tmp2194;
    wire const2430_0;
    wire[247:0] tmp2844;
    wire[7:0] tmp2895;
    wire[255:0] tmp791;
    wire[255:0] tmp2786;
    wire[255:0] tmp2195;
    wire[7:0] tmp1663;
    wire[255:0] tmp821;
    wire[7:0] tmp2366;
    wire[255:0] tmp2200;
    wire[7:0] b1_w3;
    wire const2197_0;
    wire const2550_0;
    wire[247:0] tmp2198;
    wire[247:0] tmp1917;
    wire[255:0] tmp787;
    wire[127:0] input_wire_10;
    wire[255:0] tmp2199;
    wire[7:0] b2_w3;
    wire[127:0] new_10;
    wire[127:0] tmp2897;
    wire[247:0] tmp2784;
    wire[7:0] tmp2590;
    wire[247:0] tmp2013;
    wire[255:0] tmp795;
    wire[127:0] new_5;
    wire const792_0;
    wire[255:0] tmp2845;
    wire[127:0] tmp589;
    wire[127:0] tmp1140;
    wire[247:0] tmp2170;
    wire const447_0;
    wire[255:0] tmp450;
    wire[7:0] tmp2322;
    wire[7:0] b3_w31;
    wire[7:0] tmp89;
    wire const2522_0;
    wire[7:0] tmp2380;
    wire const1025_0;
    wire[7:0] tmp1141;
    wire[247:0] tmp2210;
    wire[255:0] tmp445;
    wire[7:0] tmp2141;
    wire[7:0] tmp2950;
    wire[7:0] tmp1142;
    wire[7:0] tmp1504;
    wire[7:0] tmp1980;
    wire[255:0] tmp446;
    wire[7:0] tmp2077;
    wire[7:0] tmp853;
    wire[247:0] tmp448;
    wire[255:0] tmp2778;
    wire[255:0] tmp1313;
    wire[7:0] tmp854;
    wire[255:0] tmp421;
    wire[127:0] tmp1792;
    wire[255:0] tmp2493;
    wire[247:0] tmp2551;
    wire[255:0] tmp2441;
    wire[255:0] tmp454;
    wire const451_0;
    wire[7:0] tmp1143;
    wire[247:0] tmp452;
    wire[7:0] tmp1146;
    wire[255:0] tmp453;
    wire[7:0] tmp1920;
    wire[127:0] temp_1;
    wire[255:0] tmp1383;
    wire[127:0] temp_2;
    wire[255:0] tmp1664;
    wire[127:0] temp_3;
    wire[127:0] temp_4;
    wire[127:0] temp_5;
    wire[127:0] temp_6;
    wire[7:0] c4_w31;
    wire[127:0] temp_7;
    wire const459_0;
    wire[7:0] tmp613;
    wire[255:0] tmp462;
    wire[255:0] tmp456;
    wire[255:0] tmp1542;
    wire[127:0] temp_11;
    wire const1976_0;
    wire[255:0] tmp2010;
    wire[127:0] temp_12;
    wire[7:0] tmp1747;
    wire[127:0] temp_13;
    wire[7:0] tmp239;
    wire[127:0] temp_14;
    wire[255:0] tmp1721;
    wire[127:0] temp_15;
    wire[255:0] tmp458;
    wire const1984_0;
    wire[7:0] rc4_w11;
    wire[127:0] temp_17;
    wire[247:0] tmp460;
    wire[7:0] tmp1748;
    wire[127:0] temp_19;
    wire[127:0] temp_20;
    wire[255:0] tmp1316;
    wire[255:0] tmp461;
    wire[7:0] tmp903;
    wire[7:0] tmp1154;
    wire const2851_0;
    wire[127:0] temp_23;
    wire[7:0] tmp564;
    wire[255:0] tmp466;
    wire[7:0] tmp1029;
    wire[7:0] tmp1155;
    wire[247:0] tmp464;
    wire[255:0] tmp2235;
    wire[7:0] tmp614;
    wire[127:0] temp_27;
    wire[7:0] tmp1156;
    wire[255:0] tmp1981;
    wire[255:0] tmp465;
    wire[127:0] temp_30;
    wire const1535_0;
    wire[127:0] temp_31;
    wire[7:0] tmp1158;
    wire[7:0] tmp276;
    wire[127:0] temp_33;
    wire const2875_0;
    wire[7:0] tmp1160;
    wire[255:0] tmp2848;
    wire[127:0] temp_35;
    wire[255:0] tmp540;
    wire[127:0] temp_36;
    wire[255:0] tmp2437;
    wire[7:0] tmp1163;
    wire const1254_0;
    wire[7:0] tmp1164;
    wire[255:0] tmp1666;
    wire[255:0] tmp526;
    wire[7:0] tmp16;
    wire const2205_0;
    wire[255:0] tmp1919;
    wire[255:0] tmp2208;
    wire[255:0] tmp2519;
    wire[247:0] tmp1853;
    wire[7:0] tmp1752;
    wire[255:0] tmp794;
    wire[7:0] tmp515;
    wire[7:0] tmp2899;
    wire const1318_0;
    wire[255:0] tmp1854;
    wire[7:0] tmp2368;
    wire[7:0] tmp796;
    wire[7:0] tmp2900;
    wire const2558_0;
    wire[255:0] tmp2788;
    wire const1856_0;
    wire[7:0] tmp2177;
    wire[247:0] tmp1857;
    wire[247:0] tmp2780;
    wire[247:0] tmp1319;
    wire const1667_0;
    wire const800_0;
    wire[31:0] tmp163;
    wire const391_0;
    wire[255:0] tmp2207;
    wire[31:0] xor_w23;
    wire[7:0] tmp1754;
    wire[255:0] tmp1713;
    wire[255:0] tmp2557;
    wire[7:0] b2_w27;
    wire[7:0] b3_w27;
    wire[7:0] tmp1436;
    wire[255:0] tmp799;
    wire[7:0] tmp164;
    wire[7:0] tmp2616;
    wire[247:0] tmp801;
    wire[7:0] tmp2905;
    wire[7:0] tmp616;
    wire[255:0] tmp1861;
    wire[255:0] tmp2878;
    wire[255:0] tmp2565;
    wire const2562_0;
    wire[255:0] tmp1862;
    wire[7:0] tmp90;
    wire[255:0] tmp807;
    wire[255:0] tmp1257;
    wire const804_0;
    wire[7:0] tmp1168;
    wire[7:0] tmp1147;
    wire[255:0] tmp1863;
    wire[255:0] tmp2220;
    wire[7:0] tmp2908;
    wire[255:0] tmp806;
    wire[7:0] tmp1196;
    wire[7:0] tmp2909;
    wire[7:0] tmp167;
    wire[255:0] tmp2432;
    wire const2570_0;
    wire[255:0] tmp1999;
    wire[255:0] tmp2573;
    wire[7:0] tmp2617;
    wire[255:0] tmp2567;
    wire[7:0] tmp165;
    wire[7:0] tmp2911;
    wire[7:0] tmp2376;
    wire[255:0] tmp815;
    wire[255:0] tmp2219;
    wire[255:0] tmp422;
    wire[7:0] tmp17;
    wire[7:0] tmp2912;
    wire[7:0] rc1_w23;
    wire[7:0] tmp1144;
    wire[255:0] tmp2790;
    wire[7:0] tmp1872;
    wire const2221_0;
    wire[7:0] tmp281;
    wire[247:0] tmp2222;
    wire[255:0] tmp811;
    wire[7:0] tmp2914;
    wire[255:0] tmp1087;
    wire[255:0] tmp2572;
    wire[127:0] tmp1759;
    wire[255:0] tmp1879;
    wire[7:0] tmp2915;
    wire const1671_0;
    wire const2815_0;
    wire[255:0] tmp2577;
    wire[255:0] tmp2872;
    wire const2574_0;
    wire[7:0] tmp1438;
    wire[247:0] tmp2575;
    wire[7:0] tmp2919;
    wire[7:0] tmp91;
    wire const816_0;
    wire[255:0] tmp2576;
    wire[7:0] tmp283;
    wire[7:0] tmp2922;
    wire[255:0] tmp2226;
    wire[7:0] tmp60;
    wire[7:0] tmp2924;
    wire[255:0] tmp2015;
    wire[255:0] tmp468;
    wire[7:0] tmp284;
    wire[255:0] tmp2504;
    wire[127:0] tmp74;
    wire[7:0] tmp1450;
    wire[255:0] tmp449;
    wire[255:0] tmp2585;
    wire[7:0] tmp2957;
    wire[255:0] tmp2579;
    wire[255:0] tmp470;
    wire[7:0] tmp1440;
    wire[127:0] temp_8;
    wire[7:0] tmp1500;
    wire[7:0] tmp904;
    wire const1864_0;
    wire[255:0] tmp2580;
    wire[127:0] tmp121;
    wire[7:0] tmp11;
    wire[255:0] tmp1570;
    wire[7:0] tmp565;
    wire[7:0] tmp1501;
    wire[247:0] tmp1034;
    wire[7:0] tmp2110;
    wire[7:0] tmp286;
    wire[247:0] tmp2583;
    wire[7:0] tmp2623;
    wire[255:0] tmp478;
    wire[7:0] c2_w3;
    wire const475_0;
    wire[247:0] tmp476;
    wire[7:0] tmp62;
    wire[255:0] tmp2818;
    wire[255:0] tmp477;
    wire const2586_0;
    wire const399_0;
    wire[247:0] tmp2587;
    wire[7:0] tmp1505;
    wire[255:0] tmp1931;
    wire[255:0] tmp2588;
    wire[255:0] tmp1323;
    wire[7:0] tmp1506;
    wire[7:0] tmp2332;
    wire[7:0] b4_w31;
    wire const483_0;
    wire[255:0] tmp2520;
    wire[255:0] tmp486;
    wire[255:0] tmp2798;
    wire[255:0] tmp480;
    wire[255:0] tmp802;
    wire[7:0] tmp1508;
    wire[7:0] tmp2369;
    wire[255:0] tmp481;
    wire[255:0] tmp396;
    wire[127:0] tmp1206;
    wire[255:0] tmp2597;
    wire[7:0] tmp1509;
    wire[31:0] tmp197;
    wire[7:0] tmp215;
    wire[255:0] tmp482;
    wire[7:0] tmp1463;
    wire[7:0] tmp2379;
    wire[255:0] tmp2592;
    wire[7:0] tmp2334;
    wire[255:0] tmp2492;
    wire[255:0] tmp2593;
    wire[7:0] tmp1200;
    wire[31:0] tmp181;
    wire[247:0] tmp2595;
    wire[255:0] tmp1324;
    wire[7:0] tmp1512;
    wire const487_0;
    wire[7:0] tmp1615;
    wire[255:0] tmp2596;
    wire[7:0] tmp1513;
    wire[127:0] tmp1761;
    wire[127:0] tmp2898;
    wire[255:0] tmp2601;
    wire[31:0] shifted_w11;
    wire const2598_0;
    wire[247:0] tmp2599;
    wire const2510_0;
    wire[7:0] tmp491;
    wire[7:0] tmp1515;
    wire[7:0] tmp642;
    wire[255:0] tmp2600;
    wire[255:0] tmp2176;
    wire[7:0] tmp1228;
    wire[7:0] tmp2021;
    wire[7:0] tmp1516;
    wire[7:0] tmp2602;
    wire[255:0] tmp996;
    wire[7:0] tmp1518;
    wire[7:0] tmp2901;
    wire[7:0] tmp1519;
    wire[255:0] tmp2453;
    wire[7:0] tmp1520;
    wire[7:0] tmp1521;
    wire[127:0] tmp310;
    wire[127:0] tmp2603;
    wire const1410_0;
    wire[7:0] tmp1523;
    wire[255:0] tmp2507;
    wire[255:0] tmp2227;
    wire[7:0] tmp2079;
    wire[7:0] tmp1525;
    wire[255:0] tmp1261;
    wire[7:0] tmp1526;
    wire[127:0] tmp294;
    wire[7:0] tmp1527;
    wire[7:0] tmp1528;
    wire[247:0] tmp520;
    wire[255:0] tmp398;
    wire[7:0] tmp1529;
    wire[31:0] tmp107;
    wire[7:0] tmp1530;
    wire[7:0] tmp1145;
    wire[7:0] rc1_w31;
    wire[7:0] tmp1172;
    wire[7:0] tmp1736;
    wire[255:0] tmp2231;
    wire[7:0] tmp2022;
    wire[127:0] tmp1173;
    wire[255:0] tmp2874;
    wire[255:0] tmp1532;
    wire const1619_0;
    wire[255:0] tmp822;
    wire[127:0] tmp20;
    wire const2233_0;
    wire[255:0] tmp1538;
    wire[255:0] tmp1533;
    wire[127:0] tmp1174;
    wire[255:0] tmp2873;
    wire[255:0] tmp1534;
    wire[247:0] tmp400;
    wire[247:0] tmp1536;
    wire[127:0] tmp1175;
    wire const2173_0;
    wire[7:0] const176_0;
    wire[127:0] temp_21;
    wire[7:0] tmp1743;
    wire[255:0] tmp1537;
    wire[255:0] tmp831;
    wire[7:0] tmp2342;
    wire[247:0] tmp428;
    wire const828_0;
    wire[127:0] tmp1176;
    wire const1559_0;
    wire[255:0] tmp2244;
    wire[247:0] tmp1540;
    wire[255:0] tmp1677;
    wire[31:0] tmp178;
    wire[31:0] w0;
    wire[7:0] tmp582;
    wire[255:0] tmp1541;
    wire[255:0] tmp1638;
    wire[7:0] tmp832;
    wire[247:0] tmp1696;
    wire[31:0] tmp179;
    wire[255:0] tmp2240;
    wire[7:0] b4_w11;
    wire[255:0] tmp2166;
    wire[247:0] tmp2242;
    wire[255:0] tmp2164;
    wire const836_0;
    wire[255:0] tmp839;
    wire[7:0] const200_0;
    wire[255:0] tmp2243;
    wire[255:0] tmp1550;
    wire[127:0] temp_24;
    wire[127:0] tmp1179;
    wire[247:0] tmp2234;
    wire[255:0] tmp2248;
    wire[255:0] tmp1859;
    wire const2245_0;
    wire[247:0] tmp2246;
    wire[255:0] tmp1665;
    wire[127:0] tmp199;
    wire[255:0] tmp835;
    wire[127:0] tmp1180;
    wire[7:0] tmp2383;
    wire[255:0] tmp1546;
    wire[7:0] a4_w31;
    wire[7:0] tmp1860;
    wire[247:0] tmp2162;
    wire[247:0] tmp1548;
    wire[255:0] tmp1320;
    wire[7:0] tmp2249;
    wire[255:0] tmp2584;
    wire[127:0] tmp1181;
    wire[255:0] tmp1549;
    wire[127:0] temp_26;
    wire[255:0] tmp843;
    wire[7:0] tmp185;
    wire[7:0] tmp1445;
    wire[255:0] tmp1554;
    wire[255:0] tmp2521;
    wire const1551_0;
    wire[255:0] tmp1557;
    wire[255:0] tmp2250;
    wire[127:0] tmp195;
    wire[255:0] tmp842;
    wire[247:0] tmp1680;
    wire[7:0] tmp186;
    wire[255:0] tmp1407;
    wire[255:0] tmp2769;
    wire[255:0] tmp2251;
    wire[127:0] tmp603;
    wire[127:0] tmp1183;
    wire[255:0] tmp2252;
    wire[255:0] tmp2143;
    wire[7:0] tmp187;
    wire[7:0] tmp2384;
    wire[127:0] tmp1771;
    wire[7:0] tmp2926;
    wire[255:0] tmp2163;
    wire[7:0] tmp2927;
    wire[7:0] tmp2494;
    wire[7:0] tmp2928;
    wire[255:0] tmp1883;
    wire[7:0] tmp2930;
    wire[127:0] temp_29;
    wire[127:0] tmp2947;
    wire[127:0] tmp2931;
    wire[255:0] tmp1882;
    wire[255:0] tmp1558;
    wire[255:0] tmp502;
    wire const499_0;
    wire[255:0] tmp1681;
    wire[7:0] tmp1884;
    wire[255:0] tmp1610;
    wire[7:0] tmp1215;
    wire[255:0] tmp501;
    wire[255:0] tmp2581;
    wire[127:0] tmp2933;
    wire[7:0] tmp626;
    wire[255:0] tmp1891;
    wire[255:0] tmp1885;
    wire[255:0] tmp2517;
    wire const1133_0;
    wire[255:0] tmp2014;
    wire[255:0] tmp2483;
    wire const2863_0;
    wire[127:0] tmp2934;
    wire const507_0;
    wire[7:0] tmp467;
    wire[255:0] tmp510;
    wire[255:0] tmp1887;
    wire[7:0] tmp1447;
    wire[127:0] tmp2935;
    wire[255:0] tmp505;
    wire[7:0] tmp1152;
    wire[255:0] tmp1686;
    wire[255:0] tmp1890;
    wire[255:0] tmp506;
    wire[31:0] tmp22;
    wire[127:0] tmp2936;
    wire[255:0] tmp2569;
    wire[255:0] tmp1895;
    wire[31:0] tmp183;
    wire[247:0] tmp1893;
    wire[7:0] tmp66;
    wire[255:0] tmp509;
    wire[127:0] tmp2937;
    wire[7:0] tmp407;
    wire[255:0] tmp1894;
    wire[255:0] tmp514;
    wire[7:0] const202_0;
    wire const511_0;
    wire[247:0] tmp512;
    wire[7:0] tmp1161;
    wire[127:0] tmp2938;
    wire[255:0] tmp1626;
    wire[255:0] tmp513;
    wire const1900_0;
    wire[127:0] tmp2939;
    wire[255:0] tmp2212;
    wire[7:0] tmp1162;
    wire[7:0] tmp1746;
    wire[255:0] tmp1897;
    wire[255:0] tmp2516;
    wire[7:0] tmp189;
    wire[247:0] tmp2523;
    wire[255:0] tmp1898;
    wire[127:0] tmp2940;
    wire[255:0] tmp522;
    wire[7:0] tmp2028;
    wire[255:0] tmp1899;
    wire[31:0] concat_w19;
    wire[247:0] tmp1901;
    wire[127:0] tmp2941;
    wire[255:0] tmp1566;
    wire[255:0] tmp1902;
    wire[255:0] tmp1685;
    wire[255:0] tmp518;
    wire[31:0] tmp128;
    wire[127:0] tmp2942;
    wire const1904_0;
    wire const1563_0;
    wire[7:0] tmp1195;
    wire[7:0] tmp2116;
    wire[7:0] tmp2686;
    wire[247:0] tmp1905;
    wire[255:0] tmp774;
    wire[127:0] tmp1184;
    wire[127:0] input_wire_9;
    wire[7:0] tmp2518;
    wire[127:0] tmp2943;
    wire[247:0] tmp2527;
    wire[31:0] shifted_w31;
    wire[247:0] tmp1564;
    wire[127:0] new_9;
    wire[7:0] tmp1908;
    wire[255:0] tmp2552;
    wire[127:0] tmp2944;
    wire[127:0] tmp2348;
    wire[7:0] b1_w31;
    wire[7:0] b2_w31;
    wire[255:0] tmp2589;
    wire[127:0] tmp1186;
    wire[255:0] tmp2175;
    wire[255:0] tmp1288;
    wire const2209_0;
    wire[255:0] tmp2718;
    wire[127:0] tmp2945;
    wire[255:0] tmp408;
    wire[7:0] tmp2606;
    wire[255:0] tmp1910;
    wire[7:0] tmp848;
    wire[255:0] tmp2202;
    wire[255:0] tmp1911;
    wire[255:0] tmp1408;
    wire[31:0] w4;
    wire[7:0] tmp2902;
    wire[7:0] tmp1451;
    wire const2438_0;
    wire[247:0] tmp1913;
    wire[255:0] tmp1565;
    wire[7:0] tmp191;
    wire[255:0] tmp2144;
    wire[255:0] tmp1914;
    wire[7:0] tmp2554;
    wire[31:0] tmp55;
    wire[7:0] tmp2948;
    wire[7:0] const25_0;
    wire[7:0] tmp2610;
    wire const1916_0;
    wire[127:0] tmp846;
    wire[7:0] tmp2949;
    wire[7:0] tmp2117;
    wire[7:0] tmp2611;
    wire[7:0] tmp2030;
    wire[255:0] tmp2877;
    wire[255:0] tmp1918;
    wire[255:0] tmp2168;
    wire[7:0] tmp2612;
    wire[7:0] c2_w31;
    wire[7:0] tmp1192;
    wire[7:0] tmp2613;
    wire[255:0] tmp2203;
    wire[255:0] tmp2814;
    wire[7:0] tmp1193;
    wire[255:0] tmp2525;
    wire[247:0] tmp484;
    wire[7:0] tmp2614;
    wire const1924_0;
    wire[7:0] tmp1567;
    wire[255:0] tmp1915;
    wire[7:0] tmp1194;
    wire[7:0] tmp2615;
    wire[255:0] tmp2752;
    wire[255:0] tmp2721;
    wire[127:0] temp_9;
    wire[127:0] tmp194;
    wire[7:0] c1_w3;
    wire[7:0] const125_0;
    wire[255:0] tmp1922;
    wire[7:0] tmp2016;
    wire[255:0] tmp2003;
    wire[7:0] tmp2955;
    wire[7:0] tmp858;
    wire[7:0] tmp2956;
    wire[7:0] tmp1456;
    wire[7:0] tmp2618;
    wire[255:0] tmp2858;
    wire[7:0] tmp2081;
    wire[255:0] tmp1926;
    wire[7:0] tmp2619;
    wire[127:0] new_state;
    wire[7:0] tmp2958;
    wire[247:0] tmp1399;
    wire[7:0] tmp1457;
    wire[7:0] tmp2608;
    wire[7:0] tmp2620;
    wire[247:0] tmp1929;
    wire[7:0] tmp2959;
    wire[7:0] tmp2621;
    wire[255:0] tmp2726;
    wire[255:0] tmp1930;
    wire[127:0] tmp2353;
    wire[7:0] tmp1201;
    wire[255:0] tmp2171;
    wire[247:0] tmp2254;
    wire[247:0] tmp1668;
    wire[7:0] rc2_w31;
    wire[7:0] rc3_w31;
    wire const2723_0;
    wire[255:0] tmp2255;
    wire[255:0] tmp1562;
    wire[7:0] tmp2395;
    wire[7:0] tmp1459;
    wire[255:0] tmp1556;
    wire[255:0] tmp2260;
    wire const1571_0;
    wire const2257_0;
    wire[247:0] tmp2258;
    wire[31:0] shifted_w27;
    wire[127:0] temp_10;
    wire[7:0] tmp1749;
    wire[255:0] tmp2259;
    wire[255:0] tmp2524;
    wire[7:0] tmp1776;
    wire[247:0] tmp1560;
    wire[127:0] tmp196;
    wire[7:0] tmp580;
    wire[127:0] tmp885;
    wire[7:0] tmp2261;
    wire[255:0] tmp803;
    wire[127:0] input_wire_6;
    wire[127:0] tmp1725;
    wire[255:0] tmp1561;
    wire[7:0] tmp1461;
    wire[255:0] tmp2435;
    wire[7:0] tmp569;
    wire[31:0] tmp208;
    wire const2265_0;
    wire[255:0] tmp2268;
    wire[7:0] tmp2033;
    wire[255:0] tmp2785;
    wire[255:0] tmp2262;
    wire[127:0] tmp1772;
    wire[247:0] tmp1704;
    wire[7:0] tmp1531;
    wire[7:0] tmp820;
    wire[255:0] tmp2263;
    wire[255:0] tmp2272;
    wire[255:0] tmp2725;
    wire[255:0] tmp2264;
    wire[31:0] tmp205;
    wire[247:0] tmp2174;
    wire[247:0] tmp2266;
    wire[255:0] tmp2528;
    wire[31:0] tmp206;
    wire[7:0] a1_w35;
    wire[255:0] tmp2267;
    wire[7:0] tmp1812;
    wire[255:0] tmp1574;
    wire[255:0] tmp1568;
    wire[7:0] tmp1464;
    wire[255:0] tmp2469;
    wire const2269_0;
    wire[255:0] tmp1569;
    wire[247:0] tmp2270;
    wire[7:0] a3_w35;
    wire[255:0] tmp1289;
    wire[255:0] tmp798;
    wire[7:0] tmp1750;
    wire[255:0] tmp2271;
    wire[7:0] tmp1465;
    wire const1547_0;
    wire[247:0] tmp1572;
    wire[7:0] tmp2273;
    wire[255:0] tmp485;
    wire[7:0] tmp2727;
    wire[7:0] tmp210;
    wire[31:0] w7;
    wire[7:0] tmp2372;
    wire[127:0] tmp1482;
    wire[7:0] const77_0;
    wire[255:0] tmp1578;
    wire[7:0] tmp618;
    wire const1575_0;
    wire[7:0] tmp211;
    wire[247:0] tmp2559;
    wire[7:0] tmp2847;
    wire[127:0] tmp1466;
    wire[255:0] tmp1577;
    wire[247:0] tmp1576;
    wire[7:0] a4_w19;
    wire[7:0] tmp209;
    wire[7:0] tmp212;
    wire[7:0] tmp1579;
    wire[255:0] tmp2239;
    wire[255:0] tmp365;
    wire[255:0] tmp2882;
    wire[255:0] tmp2159;
    wire const2466_0;
    wire[31:0] shifted_w35;
    wire[255:0] tmp2279;
    wire[255:0] tmp1586;
    wire[7:0] c3_w3;
    wire[7:0] tmp2622;
    wire[7:0] tmp2397;
    wire[7:0] c4_w3;
    wire[7:0] tmp2624;
    wire[7:0] tmp864;
    wire[255:0] tmp1256;
    wire[7:0] tmp2626;
    wire[255:0] tmp2753;
    wire[255:0] tmp2211;
    wire[7:0] tmp1203;
    wire[7:0] tmp2628;
    wire[255:0] tmp739;
    wire const1001_0;
    wire[7:0] tmp2629;
    wire[7:0] tmp2630;
    wire[7:0] tmp2631;
    wire[7:0] tmp1220;
    wire[7:0] tmp2632;
    wire[255:0] tmp1867;
    wire[7:0] tmp1751;
    wire[7:0] tmp2633;
    wire[7:0] tmp2324;
    wire[7:0] tmp527;
    wire[7:0] tmp2664;
    wire[7:0] tmp2635;
    wire[255:0] tmp1617;
    wire[7:0] tmp2636;
    wire[7:0] tmp2082;
    wire[7:0] tmp2637;
    wire[7:0] tmp877;
    wire[7:0] tmp2037;
    wire[127:0] tmp2638;
    wire[7:0] tmp859;
    wire[7:0] tmp1207;
    wire[255:0] tmp1090;
    wire[255:0] tmp528;
    wire[255:0] tmp2495;
    wire[127:0] tmp880;
    wire[7:0] tmp1148;
    wire[7:0] tmp1208;
    wire[255:0] tmp529;
    wire[247:0] tmp777;
    wire[7:0] tmp1437;
    wire[7:0] tmp1209;
    wire[255:0] tmp530;
    wire[255:0] tmp1669;
    wire[7:0] tmp1210;
    wire[7:0] tmp2906;
    wire[7:0] tmp1211;
    wire[7:0] tmp2398;
    wire[255:0] tmp550;
    wire[127:0] tmp2641;
    wire[255:0] tmp538;
    wire const535_0;
    wire[247:0] tmp2563;
    wire[247:0] tmp536;
    wire[7:0] tmp1213;
    wire[31:0] substituted_w3;
    wire[255:0] tmp742;
    wire[247:0] tmp1002;
    wire[255:0] tmp1544;
    wire[255:0] tmp537;
    wire const2277_0;
    wire[7:0] tmp1214;
    wire[127:0] tmp884;
    wire[255:0] tmp2729;
    wire[127:0] new_6;
    wire[7:0] tmp539;
    wire[247:0] tmp1411;
    wire[127:0] tmp2643;
    wire[255:0] tmp1260;
    wire[255:0] tmp2436;
    wire[7:0] tmp570;
    wire[255:0] tmp2280;
    wire[7:0] tmp1216;
    wire[255:0] tmp2147;
    wire const543_0;
    wire[7:0] tmp2907;
    wire[7:0] tmp2787;
    wire[255:0] tmp546;
    wire[7:0] tmp1217;
    wire[255:0] tmp429;
    wire[7:0] tmp2951;
    wire[127:0] tmp886;
    wire[7:0] const151_0;
    wire[7:0] tmp1218;
    wire[7:0] tmp1197;
    wire[127:0] tmp2645;
    wire[255:0] tmp2564;
    wire[7:0] tmp1219;
    wire[247:0] tmp500;
    wire[255:0] tmp1092;
    wire[127:0] tmp887;
    wire[31:0] substituted_w15;
    wire[247:0] tmp544;
    wire[127:0] tmp2646;
    wire[7:0] tmp166;
    wire[255:0] tmp545;
    wire[255:0] tmp2817;
    wire[127:0] tmp888;
    wire[7:0] tmp1262;
    wire[7:0] tmp192;
    wire[7:0] tmp555;
    wire[127:0] tmp2647;
    wire[7:0] c1_w27;
    wire[7:0] tmp1222;
    wire[247:0] tmp1865;
    wire[255:0] tmp2284;
    wire const2281_0;
    wire[127:0] tmp18;
    wire[247:0] tmp745;
    wire[247:0] tmp2282;
    wire[7:0] tmp1224;
    wire[127:0] tmp2017;
    wire[255:0] tmp2275;
    wire[7:0] tmp1225;
    wire[7:0] c2_w35;
    wire[7:0] tmp1226;
    wire[7:0] tmp2566;
    wire[7:0] tmp1227;
    wire[7:0] tmp2963;
    wire[7:0] tmp2373;
    wire[255:0] tmp1127;
    wire[7:0] tmp2285;
    wire[31:0] concat_w11;
    wire[7:0] tmp1230;
    wire[7:0] tmp619;
    wire[7:0] tmp1231;
    wire[7:0] tmp1232;
    wire[7:0] tmp2047;
    wire[7:0] tmp1233;
    wire[127:0] tmp2650;
    wire[255:0] tmp2292;
    wire const519_0;
    wire[255:0] tmp2286;
    wire[7:0] tmp1237;
    wire[255:0] tmp1714;
    wire[127:0] new_11;
    wire[255:0] tmp1866;
    wire[255:0] tmp2287;
    wire[255:0] tmp1245;
    wire[255:0] tmp1095;
    wire[255:0] tmp1239;
    wire[127:0] tmp2966;
    wire[255:0] tmp2276;
    wire[7:0] b1_w35;
    wire[247:0] tmp2290;
    wire[247:0] tmp974;
    wire[247:0] tmp837;
    wire[7:0] c1_w35;
    wire const1266_0;
    wire[255:0] tmp1241;
    wire[255:0] tmp1983;
    wire[7:0] c3_w35;
    wire[7:0] tmp2039;
    wire[127:0] tmp2653;
    wire[127:0] tmp2644;
    wire[255:0] tmp2296;
    wire[7:0] tmp2213;
    wire const2293_0;
    wire[247:0] tmp2294;
    wire[7:0] tmp1442;
    wire[247:0] tmp2278;
    wire[255:0] tmp2295;
    wire[7:0] tmp1221;
    wire const1246_0;
    wire[7:0] tmp2910;
    wire[7:0] tmp2655;
    wire[7:0] tmp2297;
    wire[7:0] tmp748;
    wire[7:0] tmp1510;
    wire[7:0] tmp2073;
    wire[7:0] tmp2656;
    wire const1703_0;
    wire[127:0] tmp220;
    wire[255:0] tmp2738;
    wire[127:0] tmp2605;
    wire const2301_0;
    wire[7:0] tmp860;
    wire[255:0] tmp2304;
    wire[255:0] tmp1990;
    wire[255:0] tmp2298;
    wire[255:0] tmp2496;
    wire[7:0] tmp2658;
    wire[7:0] tmp1149;
    wire[255:0] tmp2299;
    wire const2735_0;
    wire[7:0] tmp2659;
    wire[255:0] tmp1251;
    wire[127:0] tmp1767;
    wire[31:0] shifted_w23;
    wire[255:0] tmp2300;
    wire[7:0] tmp2660;
    wire[31:0] tmp213;
    wire[247:0] tmp2302;
    wire[7:0] b2_w35;
    wire const812_0;
    wire[7:0] tmp2661;
    wire[255:0] tmp1253;
    wire[7:0] tmp2401;
    wire[7:0] rc2_w35;
    wire[255:0] tmp433;
    wire[247:0] tmp1255;
    wire[7:0] tmp2040;
    wire[255:0] tmp2308;
    wire[7:0] const223_9;
    wire[255:0] tmp1292;
    wire[7:0] c2_w27;
    wire[7:0] tmp2663;
    wire const2803_0;
    wire[127:0] tmp224;
    wire const547_0;
    wire[247:0] tmp548;
    wire const2731_0;
    wire[255:0] tmp1870;
    wire[7:0] tmp290;
    wire[255:0] tmp1581;
    wire[255:0] tmp1412;
    wire[255:0] tmp549;
    wire const752_0;
    wire[7:0] tmp1896;
    wire const1936_0;
    wire[7:0] tmp863;
    wire[255:0] tmp1706;
    wire[255:0] tmp1939;
    wire[255:0] tmp1933;
    wire[7:0] tmp2023;
    wire[7:0] c4_w27;
    wire[247:0] tmp1833;
    wire[255:0] tmp1265;
    wire[7:0] tmp2952;
    wire[255:0] tmp1934;
    wire[127:0] tmp552;
    wire[7:0] const152_0;
    wire[7:0] tmp1198;
    wire[255:0] tmp1935;
    wire[31:0] substituted_w27;
    wire const1587_0;
    wire[247:0] tmp1937;
    wire[7:0] b1_w23;
    wire[255:0] tmp1325;
    wire[7:0] tmp1202;
    wire[255:0] tmp1938;
    wire[7:0] tmp2903;
    wire[7:0] b3_w35;
    wire[127:0] tmp553;
    wire[255:0] tmp2224;
    wire[255:0] tmp2822;
    wire[255:0] tmp1943;
    wire[7:0] b2_w23;
    wire const1940_0;
    wire[247:0] tmp1941;
    wire[7:0] tmp2041;
    wire[7:0] tmp2739;
    wire const1595_0;
    wire[7:0] tmp2341;
    wire[255:0] tmp2850;
    wire[255:0] tmp1598;
    wire[255:0] tmp1592;
    wire const2161_0;
    wire[255:0] tmp1580;
    wire[7:0] tmp1944;
    wire[127:0] input_wire_2;
    wire[7:0] tmp865;
    wire[255:0] tmp1593;
    wire[247:0] tmp2571;
    wire[7:0] tmp1483;
    wire[127:0] tmp1470;
    wire[7:0] b4_w23;
    wire[255:0] tmp457;
    wire[255:0] tmp1594;
    wire[255:0] tmp2508;
    wire[255:0] tmp1951;
    wire[7:0] tmp572;
    wire[255:0] tmp1393;
    wire[127:0] tmp620;
    wire[255:0] tmp1945;
    wire[7:0] tmp558;
    wire[255:0] tmp2183;
    wire[255:0] tmp1946;
    wire[255:0] tmp1993;
    wire[7:0] tmp559;
    wire[7:0] tmp334;
    wire[255:0] tmp1947;
    wire[255:0] tmp1927;
    wire const1599_0;
    wire[127:0] tmp2054;
    wire[247:0] tmp1949;
    wire[255:0] tmp2303;
    wire[7:0] tmp561;
    wire[255:0] tmp2555;
    wire[31:0] tmp133;
    wire[255:0] tmp1950;
    wire[247:0] tmp1391;
    wire[7:0] b4_w35;
    wire[7:0] tmp562;
    wire const1876_0;
    wire[255:0] tmp1955;
    wire const1952_0;
    wire[7:0] tmp808;
    wire const1105_0;
    wire[247:0] tmp1953;
    wire[255:0] tmp2238;
    wire[7:0] tmp869;
    wire const1607_0;
    wire const2743_0;
    wire[127:0] temp_18;
    wire[247:0] tmp1415;
    wire[255:0] tmp1604;
    wire[7:0] tmp912;
    wire[255:0] tmp1108;
    wire[7:0] tmp1956;
    wire[127:0] tmp2310;
    wire[7:0] tmp335;
    wire[255:0] tmp1605;
    wire[255:0] tmp2151;
    wire[7:0] tmp566;
    wire[255:0] tmp1873;
    wire[127:0] temp_39;
    wire[255:0] tmp1102;
    wire const1960_0;
    wire[127:0] tmp889;
    wire[7:0] tmp573;
    wire[7:0] tmp871;
    wire[255:0] tmp1957;
    wire[7:0] tmp2309;
    wire[255:0] tmp1263;
    wire[7:0] tmp2916;
    wire[31:0] w3;
    wire[7:0] tmp861;
    wire[255:0] tmp1958;
    wire[247:0] tmp1271;
    wire[127:0] tmp890;
    wire[255:0] tmp2497;
    wire[31:0] w6;
    wire[7:0] tmp872;
    wire[7:0] tmp1150;
    wire[255:0] tmp1959;
    wire[31:0] tmp5;
    wire[7:0] tmp2693;
    wire[7:0] tmp2917;
    wire const1326_0;
    wire[247:0] tmp1961;
    wire[31:0] tmp7;
    wire[127:0] tmp895;
    wire[127:0] input_wire_8;
    wire[255:0] tmp1962;
    wire[255:0] tmp2452;
    wire[7:0] tmp214;
    wire[127:0] new_8;
    wire[7:0] tmp2918;
    wire[127:0] tmp2311;
    wire[247:0] tmp2820;
    wire const1964_0;
    wire[255:0] tmp1103;
    wire[7:0] tmp2404;
    wire[247:0] tmp1965;
    wire[7:0] tmp2470;
    wire const1069_0;
    wire[127:0] tmp2312;
    wire[7:0] tmp874;
    wire[7:0] a1_w3;
    wire[255:0] tmp1966;
    wire[255:0] tmp1297;
    wire[7:0] a3_w3;
    wire[7:0] a4_w3;
    wire[127:0] tmp19;
    wire[247:0] tmp1997;
    wire[7:0] tmp1968;
    wire[7:0] tmp2313;
    wire[31:0] xor_w19;
    wire[7:0] tmp875;
    wire[31:0] tmp233;
    wire[31:0] xor_w31;
    wire[7:0] tmp2920;
    wire[7:0] tmp2314;
    wire[7:0] tmp10;
    wire[255:0] tmp1975;
    wire[255:0] tmp1969;
    wire[255:0] tmp1640;
    wire[7:0] tmp337;
    wire[7:0] tmp234;
    wire[7:0] tmp2921;
    wire[7:0] tmp2316;
    wire[255:0] tmp1834;
    wire[255:0] tmp759;
    wire[7:0] tmp2953;
    wire[255:0] tmp1035;
    wire[7:0] tmp2317;
    wire[127:0] tmp2654;
    wire[31:0] concat_w23;
    wire[7:0] tmp1199;
    wire[7:0] tmp2095;
    wire[247:0] tmp1973;
    wire[255:0] tmp2742;
    wire[255:0] tmp1329;
    wire[7:0] tmp2318;
    wire[7:0] tmp1799;
    wire[127:0] tmp2355;
    wire[255:0] tmp1998;
    wire[255:0] tmp1974;
    wire[7:0] tmp2319;
    wire[247:0] tmp2455;
    wire[31:0] shifted_w3;
    wire[7:0] tmp899;
    wire[7:0] tmp2923;
    wire[7:0] tmp2320;
    wire[255:0] tmp2160;
    wire[247:0] tmp757;
    wire[7:0] tmp900;
    wire[255:0] tmp489;
    wire[7:0] tmp1322;
    wire[7:0] tmp2321;
    wire[7:0] tmp338;
    wire[255:0] tmp1978;
    wire[7:0] b3_w3;
    wire[255:0] tmp2757;
    wire[7:0] b4_w3;
    wire[127:0] tmp1775;
    wire[7:0] tmp14;
    wire[7:0] tmp902;
    wire[255:0] tmp1923;
    wire const1691_0;
    wire[255:0] tmp521;
    wire[7:0] tmp2323;
    wire[127:0] tmp896;
    wire[7:0] b1_w39;
    wire[7:0] tmp2925;
    wire[7:0] tmp15;
    wire[255:0] tmp1987;
    wire[7:0] tmp623;
    wire[7:0] tmp2375;
    wire[7:0] b4_w39;
    wire[255:0] tmp2500;
    wire[7:0] tmp2325;
    wire[7:0] tmp575;
    wire[255:0] tmp2456;
    wire[255:0] tmp1701;
    wire[7:0] tmp1797;
    wire[255:0] tmp1606;
    wire[127:0] tmp1774;
    wire[7:0] tmp2326;
    wire[255:0] tmp1107;
    wire[247:0] tmp1608;
    wire[247:0] tmp2499;
    wire[31:0] tmp153;
    wire[7:0] tmp568;
    wire[255:0] tmp1609;
    wire[7:0] tmp2695;
    wire[7:0] tmp1498;
    wire[247:0] tmp781;
    wire[7:0] tmp2328;
    wire const1278_0;
    wire[127:0] tmp2649;
    wire[255:0] tmp1614;
    wire[7:0] tmp560;
    wire[255:0] tmp2531;
    wire[127:0] tmp2639;
    wire[255:0] tmp1673;
    wire[7:0] tmp2329;
    wire[7:0] tmp2330;
    wire[255:0] tmp2745;
    wire[7:0] tmp2331;
    wire[255:0] tmp1613;
    wire[255:0] tmp1281;
    wire[7:0] tmp2406;
    wire[7:0] tmp2333;
    wire[255:0] tmp2765;
    wire[255:0] tmp1066;
    wire[7:0] tmp2458;
    wire const2594_0;
    wire[7:0] tmp2335;
    wire[255:0] tmp2132;
    wire[7:0] tmp2336;
    wire[247:0] tmp1295;
    wire[7:0] tmp2337;
    wire[255:0] tmp1416;
    wire[7:0] tmp2338;
    wire[7:0] tmp760;
    wire[7:0] tmp2339;
    wire[7:0] tmp2340;
    wire[127:0] new_7;
    wire[255:0] tmp1622;
    wire const2767_0;
    wire[7:0] tmp2153;
    wire[255:0] tmp1616;
    wire const2582_0;
    wire const1840_0;
    wire[7:0] tmp2343;
    wire[7:0] tmp2344;
    wire[127:0] tmp2361;
    wire[255:0] tmp1963;
    wire[127:0] tmp2345;
    wire[7:0] tmp576;
    wire[127:0] tmp881;
    wire[7:0] tmp621;
    wire[7:0] tmp1153;
    wire[255:0] tmp1618;
    wire[31:0] tmp229;
    wire[7:0] tmp2389;
    wire[127:0] tmp21;
    wire[7:0] tmp862;
    wire[247:0] tmp1620;
    wire[7:0] c1_w23;
    wire const435_0;
    wire[127:0] tmp2346;
    wire[247:0] tmp1612;
    wire[255:0] tmp1397;
    wire[7:0] tmp1151;
    wire[255:0] tmp1621;
    wire[127:0] tmp588;
    wire[7:0] tmp2627;
    wire[127:0] tmp2347;
    wire const1623_0;
    wire[247:0] tmp1624;
    wire[127:0] tmp2640;
    wire[7:0] rc1_w3;
    wire[7:0] tmp2662;
    wire[7:0] rc2_w3;
    wire[255:0] tmp1625;
    wire[255:0] tmp2821;
    wire[7:0] rc4_w3;
    wire[7:0] const23_1;
    wire[7:0] tmp1627;
    wire const2462_0;
    wire[127:0] tmp24;
    wire[255:0] tmp655;
    wire[127:0] tmp2349;
    wire[7:0] tmp2390;
    wire[255:0] tmp2214;
    wire[127:0] temp_22;
    wire[255:0] tmp2247;
    wire[255:0] tmp1111;
    wire const1631_0;
    wire[247:0] tmp1925;
    wire[7:0] tmp2078;
    wire[7:0] rc3_w19;
    wire[127:0] tmp2350;
    wire[7:0] tmp855;
    wire[7:0] const26_0;
    wire[7:0] tmp1651;
    wire[247:0] tmp472;
    wire const2145_0;
    wire[7:0] tmp2609;
    wire[7:0] tmp2913;
    wire[7:0] tmp2327;
    wire[255:0] tmp1629;
    wire[127:0] tmp1471;
    wire[7:0] const27_0;
    wire[127:0] tmp2351;
    wire[7:0] tmp577;
    wire[7:0] tmp342;
    wire[255:0] tmp1630;
    wire[31:0] concat_w3;
    wire[247:0] tmp990;
    wire[247:0] tmp1632;
    wire[255:0] tmp2307;
    wire[127:0] tmp143;
    wire[7:0] tmp2954;
    wire const2486_0;
    wire const1583_0;
    wire[7:0] tmp111;
    wire[255:0] tmp1400;
    wire[255:0] tmp1982;
    wire[255:0] tmp2123;
    wire[255:0] tmp1921;
    wire const1258_0;
    wire[7:0] tmp2391;
    wire[247:0] tmp1259;
    wire[247:0] tmp2306;
    wire[7:0] tmp2665;
    wire[247:0] tmp1279;
    wire[247:0] tmp1985;
    wire[7:0] tmp2666;
    wire[255:0] tmp473;
    wire[255:0] tmp1986;
    wire[247:0] tmp841;
    wire[7:0] tmp2667;
    wire[7:0] tmp2408;
    wire[255:0] tmp2560;
    wire[255:0] tmp1991;
    wire[255:0] tmp2460;
    wire[255:0] tmp2591;
    wire[7:0] tmp2668;
    wire[247:0] tmp1989;
    wire[255:0] tmp991;
    wire[255:0] tmp2762;
    wire[255:0] tmp1269;
    wire[7:0] tmp2669;
    wire[255:0] tmp2011;
    wire[7:0] b3_w11;
    wire[255:0] tmp1582;
    wire[255:0] tmp1405;
    wire[7:0] tmp2670;
    wire[7:0] tmp1992;
    wire[7:0] tmp2392;
    wire[255:0] tmp810;
    wire[7:0] tmp1727;
    wire[127:0] tmp2671;
    wire[255:0] tmp2005;
    wire[247:0] tmp1869;
    wire[255:0] tmp2505;
    wire[247:0] tmp1267;
    wire[7:0] tmp578;
    wire[127:0] tmp883;
    wire const1996_0;
    wire[7:0] tmp2672;
    wire[255:0] tmp2411;
    wire[255:0] tmp2789;
    wire[7:0] tmp2673;
    wire const1037_0;
    wire[255:0] tmp1994;
    wire[255:0] tmp2461;
    wire[127:0] tmp847;
    wire const1270_0;
    wire[7:0] tmp2674;
    wire[255:0] tmp1690;
    wire[247:0] tmp2756;
    wire[255:0] tmp1995;
    wire[7:0] tmp2904;
    wire const1117_0;
    wire[7:0] tmp2675;
    wire[255:0] tmp2532;
    wire[127:0] tmp2642;
    wire[7:0] tmp1675;
    wire[7:0] tmp2676;
    wire[7:0] tmp2393;
    wire[255:0] tmp1670;
    wire[255:0] tmp2006;
    wire[7:0] tmp2409;
    wire[7:0] tmp2677;
    wire const2474_0;
    wire const2000_0;
    wire[247:0] tmp2463;
    wire[247:0] tmp2001;
    wire[127:0] tmp169;
    wire[7:0] tmp2678;
    wire[255:0] tmp1296;
    wire const2759_0;
    wire[255:0] tmp1275;
    wire[255:0] tmp2002;
    wire[247:0] tmp817;
    wire[7:0] rc2_w27;
    wire[255:0] tmp525;
    wire[7:0] tmp2679;
    wire[255:0] tmp2761;
    wire const523_0;
    wire[255:0] tmp1276;
    wire[255:0] tmp1404;
    wire[7:0] tmp2004;
    wire[7:0] c4_w35;
    wire[7:0] rc4_w31;
    wire[7:0] tmp2680;
    wire[255:0] tmp2730;
    wire[255:0] tmp1277;
    wire[7:0] const173_7;
    wire[7:0] tmp2681;
    wire[255:0] tmp2445;
    wire const2502_0;
    wire const2008_0;
    wire[7:0] tmp579;
    wire[7:0] tmp348;
    wire[7:0] tmp622;
    wire[247:0] tmp2892;
    wire[7:0] tmp2682;
    wire[255:0] tmp1835;
    wire[7:0] tmp2394;
    wire[255:0] tmp2556;
    wire[255:0] tmp2007;
    wire[7:0] tmp2683;
    wire[247:0] tmp1038;
    wire[7:0] tmp1932;
    wire const1282_0;
    wire[255:0] tmp2464;
    wire[7:0] tmp1229;
    wire[247:0] tmp1283;
    wire[7:0] tmp2684;
    wire[255:0] tmp1693;

    reg[255:0] mem_4[255:0];
    reg[255:0] mem_3[255:0];
    reg[127:0] mem_2[255:0];
    reg[127:0] mem_1[255:0];

    assign const126_0 = 0;
    assign const1338_0 = 0;
    assign const2887_0 = 0;
    assign const1539_0 = 0;
    assign const427_0 = 0;
    assign const1414_0 = 0;
    assign const252_0 = 0;
    assign const1571_0 = 0;
    assign const2546_0 = 0;
    assign const2731_0 = 0;
    assign const2125_0 = 0;
    assign const1254_0 = 0;
    assign const2426_0 = 0;
    assign const2430_0 = 0;
    assign const1635_0 = 0;
    assign const2197_0 = 0;
    assign const1928_0 = 0;
    assign const1270_0 = 0;
    assign const1936_0 = 0;
    assign const2771_0 = 0;
    assign const2193_0 = 0;
    assign const1924_0 = 0;
    assign const2145_0 = 0;
    assign const2558_0 = 0;
    assign const423_0 = 0;
    assign const732_0 = 0;
    assign const2879_0 = 0;
    assign const2851_0 = 0;
    assign const1258_0 = 0;
    assign const2723_0 = 0;
    assign const2185_0 = 0;
    assign const2478_0 = 0;
    assign const1916_0 = 0;
    assign const2233_0 = 0;
    assign const2209_0 = 0;
    assign const2526_0 = 0;
    assign const459_0 = 0;
    assign const1422_0 = 0;
    assign const1988_0 = 0;
    assign const2205_0 = 0;
    assign const2855_0 = 0;
    assign const1832_0 = 0;
    assign const2711_0 = 0;
    assign const2133_0 = 0;
    assign const1996_0 = 0;
    assign const198_8 = 8;
    assign const1342_0 = 0;
    assign const1940_0 = 0;
    assign const2594_0 = 0;
    assign const1643_0 = 0;
    assign const1844_0 = 0;
    assign const27_0 = 0;
    assign const1398_0 = 0;
    assign const2281_0 = 0;
    assign const1912_0 = 0;
    assign const1266_0 = 0;
    assign const2173_0 = 0;
    assign const176_0 = 0;
    assign const2707_0 = 0;
    assign const2438_0 = 0;
    assign const2169_0 = 0;
    assign const523_0 = 0;
    assign const1073_0 = 0;
    assign const2257_0 = 0;
    assign const672_0 = 0;
    assign const828_0 = 0;
    assign const2767_0 = 0;
    assign const2241_0 = 0;
    assign const2229_0 = 0;
    assign const1013_0 = 0;
    assign const1840_0 = 0;
    assign const973_0 = 0;
    assign const1575_0 = 0;
    assign const125_0 = 0;
    assign const1109_0 = 0;
    assign const1049_0 = 0;
    assign const2217_0 = 0;
    assign const1350_0 = 0;
    assign const2562_0 = 0;
    assign const2783_0 = 0;
    assign const2161_0 = 0;
    assign const1426_0 = 0;
    assign const768_0 = 0;
    assign const439_0 = 0;
    assign const127_0 = 0;
    assign const2137_0 = 0;
    assign const953_0 = 0;
    assign const435_0 = 0;
    assign const780_0 = 0;
    assign const2843_0 = 0;
    assign const543_0 = 0;
    assign const1647_0 = 0;
    assign const728_0 = 0;
    assign const152_0 = 0;
    assign const836_0 = 0;
    assign const2574_0 = 0;
    assign const2181_0 = 0;
    assign const2570_0 = 0;
    assign const1559_0 = 0;
    assign const447_0 = 0;
    assign const2891_0 = 0;
    assign const708_0 = 0;
    assign const2735_0 = 0;
    assign const471_0 = 0;
    assign const2490_0 = 0;
    assign const2586_0 = 0;
    assign const1595_0 = 0;
    assign const2791_0 = 0;
    assign const977_0 = 0;
    assign const1390_0 = 0;
    assign const2867_0 = 0;
    assign const1659_0 = 0;
    assign const1033_0 = 0;
    assign const2598_0 = 0;
    assign const1354_0 = 0;
    assign const200_0 = 0;
    assign const1655_0 = 0;
    assign const2462_0 = 0;
    assign const387_0 = 0;
    assign const684_0 = 0;
    assign const1607_0 = 0;
    assign const23_1 = 1;
    assign const2305_0 = 0;
    assign const463_0 = 0;
    assign const1876_0 = 0;
    assign const175_0 = 0;
    assign const2442_0 = 0;
    assign const1892_0 = 0;
    assign const1085_0 = 0;
    assign const2819_0 = 0;
    assign const2221_0 = 0;
    assign const363_0 = 0;
    assign const1888_0 = 0;
    assign const1105_0 = 0;
    assign const2815_0 = 0;
    assign const2253_0 = 0;
    assign const985_0 = 0;
    assign const1619_0 = 0;
    assign const989_0 = 0;
    assign const2875_0 = 0;
    assign const26_0 = 0;
    assign const692_0 = 0;
    assign const2719_0 = 0;
    assign const1631_0 = 0;
    assign const1362_0 = 0;
    assign const2277_0 = 0;
    assign const2450_0 = 0;
    assign const2795_0 = 0;
    assign const2831_0 = 0;
    assign const949_0 = 0;
    assign const415_0 = 0;
    assign const2121_0 = 0;
    assign const1852_0 = 0;
    assign const1828_0 = 0;
    assign const227_0 = 0;
    assign const2149_0 = 0;
    assign const2008_0 = 0;
    assign const251_0 = 0;
    assign const744_0 = 0;
    assign const840_0 = 0;
    assign const2293_0 = 0;
    assign const812_0 = 0;
    assign const2486_0 = 0;
    assign const1583_0 = 0;
    assign const1093_0 = 0;
    assign const2839_0 = 0;
    assign const1960_0 = 0;
    assign const1117_0 = 0;
    assign const2827_0 = 0;
    assign const150_0 = 0;
    assign const1045_0 = 0;
    assign const1868_0 = 0;
    assign const2582_0 = 0;
    assign const1314_0 = 0;
    assign const1864_0 = 0;
    assign const248_10 = 10;
    assign const1535_0 = 0;
    assign const2747_0 = 0;
    assign const2522_0 = 0;
    assign const824_0 = 0;
    assign const226_0 = 0;
    assign const403_0 = 0;
    assign const668_0 = 0;
    assign const2012_0 = 0;
    assign const2466_0 = 0;
    assign const800_0 = 0;
    assign const1611_0 = 0;
    assign const1290_0 = 0;
    assign const499_0 = 0;
    assign const1410_0 = 0;
    assign const250_0 = 0;
    assign const1326_0 = 0;
    assign const1366_0 = 0;
    assign const752_0 = 0;
    assign const1984_0 = 0;
    assign const1880_0 = 0;
    assign const1667_0 = 0;
    assign const2807_0 = 0;
    assign const2534_0 = 0;
    assign const2289_0 = 0;
    assign const2779_0 = 0;
    assign const1948_0 = 0;
    assign const475_0 = 0;
    assign const519_0 = 0;
    assign const177_0 = 0;
    assign const1599_0 = 0;
    assign const1121_0 = 0;
    assign const51_0 = 0;
    assign const2269_0 = 0;
    assign const411_0 = 0;
    assign const148_6 = 6;
    assign const2265_0 = 0;
    assign const1081_0 = 0;
    assign const1719_0 = 0;
    assign const1133_0 = 0;
    assign const1069_0 = 0;
    assign const997_0 = 0;
    assign const1679_0 = 0;
    assign const965_0 = 0;
    assign const2863_0 = 0;
    assign const1318_0 = 0;
    assign const507_0 = 0;
    assign const1061_0 = 0;
    assign const535_0 = 0;
    assign const1374_0 = 0;
    assign const2498_0 = 0;
    assign const1242_0 = 0;
    assign const1695_0 = 0;
    assign const531_0 = 0;
    assign const1402_0 = 0;
    assign const379_0 = 0;
    assign const2157_0 = 0;
    assign const2245_0 = 0;
    assign const1294_0 = 0;
    assign const2474_0 = 0;
    assign const720_0 = 0;
    assign const1129_0 = 0;
    assign const151_0 = 0;
    assign const1306_0 = 0;
    assign const1856_0 = 0;
    assign const816_0 = 0;
    assign const2514_0 = 0;
    assign const1671_0 = 0;
    assign const547_0 = 0;
    assign const2538_0 = 0;
    assign const2510_0 = 0;
    assign const680_0 = 0;
    assign const704_0 = 0;
    assign const391_0 = 0;
    assign const98_4 = 4;
    assign const1587_0 = 0;
    assign const1021_0 = 0;
    assign const100_0 = 0;
    assign const764_0 = 0;
    assign const2759_0 = 0;
    assign const1278_0 = 0;
    assign const52_0 = 0;
    assign const1976_0 = 0;
    assign const1246_0 = 0;
    assign const1972_0 = 0;
    assign const1001_0 = 0;
    assign const2414_0 = 0;
    assign const2454_0 = 0;
    assign const73_3 = 3;
    assign const1551_0 = 0;
    assign const75_0 = 0;
    assign const2550_0 = 0;
    assign const1547_0 = 0;
    assign const656_0 = 0;
    assign const2743_0 = 0;
    assign const511_0 = 0;
    assign const2000_0 = 0;
    assign const776_0 = 0;
    assign const1302_0 = 0;
    assign const1057_0 = 0;
    assign const2301_0 = 0;
    assign const483_0 = 0;
    assign const102_0 = 0;
    assign const1097_0 = 0;
    assign const1900_0 = 0;
    assign const1282_0 = 0;
    assign const48_2 = 2;
    assign const2755_0 = 0;
    assign const223_9 = 9;
    assign const50_0 = 0;
    assign const1715_0 = 0;
    assign const76_0 = 0;
    assign const1563_0 = 0;
    assign const123_5 = 5;
    assign const1009_0 = 0;
    assign const804_0 = 0;
    assign const367_0 = 0;
    assign const1330_0 = 0;
    assign const375_0 = 0;
    assign const77_0 = 0;
    assign const740_0 = 0;
    assign const25_0 = 0;
    assign const1386_0 = 0;
    assign const173_7 = 7;
    assign const1037_0 = 0;
    assign const1707_0 = 0;
    assign const2502_0 = 0;
    assign const1623_0 = 0;
    assign const1378_0 = 0;
    assign const1025_0 = 0;
    assign const2418_0 = 0;
    assign const1952_0 = 0;
    assign const1691_0 = 0;
    assign const495_0 = 0;
    assign const202_0 = 0;
    assign const696_0 = 0;
    assign const756_0 = 0;
    assign const487_0 = 0;
    assign const1703_0 = 0;
    assign const1683_0 = 0;
    assign const660_0 = 0;
    assign const399_0 = 0;
    assign const792_0 = 0;
    assign const201_0 = 0;
    assign const961_0 = 0;
    assign const716_0 = 0;
    assign const1964_0 = 0;
    assign const101_0 = 0;
    assign const225_0 = 0;
    assign const788_0 = 0;
    assign const2803_0 = 0;
    assign const1904_0 = 0;
    assign const451_0 = 0;
    assign tmp2487 = {const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0, const2486_0};
    assign tmp392 = {const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0, const391_0};
        assign tmp2167 = mem_4[tmp2091];
        assign tmp2354 = mem_1[tmp2322];
    assign tmp1029 = {tmp1028[0], tmp1028[1], tmp1028[2], tmp1028[3], tmp1028[4], tmp1028[5], tmp1028[6], tmp1028[7]};
    assign b2_w7 = tmp40;
    assign tmp311 = {temp_1[120], temp_1[121], temp_1[122], temp_1[123], temp_1[124], temp_1[125], temp_1[126], temp_1[127]};
        assign tmp1850 = mem_4[tmp1796];
    assign tmp393 = {tmp392, tmp329};
    assign tmp1047 = {tmp1046, tmp924};
    assign tmp1415 = {const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0, const1414_0};
    assign tmp339 = {temp_2[32], temp_2[33], temp_2[34], temp_2[35], temp_2[36], temp_2[37], temp_2[38], temp_2[39]};
    assign tmp1797 = {temp_22[88], temp_22[89], temp_22[90], temp_22[91], temp_22[92], temp_22[93], temp_22[94], temp_22[95]};
        assign tmp1774 = mem_1[tmp1742];
        assign tmp1066 = mem_3[tmp924];
    assign tmp1262 = {tmp1261[0], tmp1261[1], tmp1261[2], tmp1261[3], tmp1261[4], tmp1261[5], tmp1261[6], tmp1261[7]};
    assign tmp400 = {const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0, const399_0};
    assign tmp1542 = tmp1538 ^ tmp1541;
    assign tmp56 = tmp55 ^ w5;
    assign tmp1162 = tmp1178;
    assign tmp2307 = {tmp2306, tmp2100};
    assign tmp2308 = tmp2304 ^ tmp2307;
    assign tmp570 = {temp_4[0], temp_4[1], temp_4[2], temp_4[3], temp_4[4], temp_4[5], temp_4[6], temp_4[7]};
    assign tmp256 = tmp255 ^ tmp231;
        assign tmp2884 = mem_3[tmp2687];
    assign tmp1632 = {const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0, const1631_0};
    assign tmp2608 = {temp_32[104], temp_32[105], temp_32[106], temp_32[107], temp_32[108], temp_32[109], temp_32[110], temp_32[111]};
        assign tmp1252 = mem_4[tmp1209];
    assign tmp462 = tmp458 ^ tmp461;
    assign tmp2721 = {tmp2720, tmp2675};
    assign tmp2434 = {tmp2433[0], tmp2433[1], tmp2433[2], tmp2433[3], tmp2433[4], tmp2433[5], tmp2433[6], tmp2433[7]};
    assign tmp1159 = tmp1175;
    assign tmp2401 = tmp2494;
        assign tmp2263 = mem_4[tmp2099];
    assign tmp1443 = {temp_16[48], temp_16[49], temp_16[50], temp_16[51], temp_16[52], temp_16[53], temp_16[54], temp_16[55]};
    assign tmp2367 = {temp_29[80], temp_29[81], temp_29[82], temp_29[83], temp_29[84], temp_29[85], temp_29[86], temp_29[87]};
    assign tmp349 = tmp431;
        assign tmp2359 = mem_1[tmp2327];
    assign tmp1859 = tmp1855 ^ tmp1858;
    assign tmp1113 = {tmp1112[0], tmp1112[1], tmp1112[2], tmp1112[3], tmp1112[4], tmp1112[5], tmp1112[6], tmp1112[7]};
    assign tmp795 = tmp791 ^ tmp794;
        assign tmp409 = mem_4[tmp333];
    assign tmp1586 = tmp1582 ^ tmp1585;
    assign tmp1975 = tmp1971 ^ tmp1974;
        assign tmp737 = mem_3[tmp628];
        assign tmp2649 = mem_1[tmp2617];
    assign tmp647 = tmp784;
    assign tmp461 = {tmp460, tmp338};
    assign tmp1805 = {temp_22[24], temp_22[25], temp_22[26], temp_22[27], temp_22[28], temp_22[29], temp_22[30], temp_22[31]};
        assign tmp373 = mem_4[tmp330];
    assign tmp1796 = {temp_22[96], temp_22[97], temp_22[98], temp_22[99], temp_22[100], temp_22[101], temp_22[102], temp_22[103]};
        assign tmp2118 = mem_3[tmp2086];
    assign tmp1747 = tmp1763;
    assign tmp988 = tmp984 ^ tmp987;
        assign tmp124 = mem_2[const123_5];
    assign tmp2114 = tmp2273;
    assign tmp1663 = {tmp1662[0], tmp1662[1], tmp1662[2], tmp1662[3], tmp1662[4], tmp1662[5], tmp1662[6], tmp1662[7]};
    assign tmp1974 = {tmp1973, tmp1807};
    assign tmp2004 = {tmp2003[0], tmp2003[1], tmp2003[2], tmp2003[3], tmp2003[4], tmp2003[5], tmp2003[6], tmp2003[7]};
    assign tmp254 = concat_w39 ^ substituted_w39;
        assign tmp1969 = mem_3[tmp1805];
    assign tmp2948 = {temp_37[120], temp_37[121], temp_37[122], temp_37[123], temp_37[124], temp_37[125], temp_37[126], temp_37[127]};
    assign tmp1145 = {temp_12[88], temp_12[89], temp_12[90], temp_12[91], temp_12[92], temp_12[93], temp_12[94], temp_12[95]};
    assign tmp2930 = tmp2946;
    assign temp_6 = tmp620;
        assign tmp1676 = mem_3[tmp1512];
    assign tmp1210 = {temp_14[96], temp_14[97], temp_14[98], temp_14[99], temp_14[100], temp_14[101], temp_14[102], temp_14[103]};
        assign tmp2752 = mem_3[tmp2676];
    assign tmp518 = tmp516 ^ tmp517;
    assign tmp158 = tmp157 ^ tmp133;
    assign tmp180 = tmp155 ^ xor_w27;
    assign tmp2528 = {tmp2527, tmp2387};
        assign tmp893 = mem_1[tmp861];
    assign tmp362 = tmp360 ^ tmp361;
        assign tmp883 = mem_1[tmp851];
        assign tmp1480 = mem_1[tmp1448];
    assign tmp2481 = tmp2477 ^ tmp2480;
    assign tmp2583 = {const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0, const2582_0};
    assign tmp1191 = {temp_13[112], temp_13[113], temp_13[114], temp_13[115], temp_13[116], temp_13[117], temp_13[118], temp_13[119]};
    assign tmp380 = {const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0, const379_0};
    assign tmp691 = tmp689 ^ tmp690;
    assign tmp2368 = {temp_29[72], temp_29[73], temp_29[74], temp_29[75], temp_29[76], temp_29[77], temp_29[78], temp_29[79]};
    assign tmp2563 = {const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0, const2562_0};
    assign tmp2902 = {temp_36[96], temp_36[97], temp_36[98], temp_36[99], temp_36[100], temp_36[101], temp_36[102], temp_36[103]};
    assign temp_4 = new_2;
    assign tmp2590 = {tmp2589[0], tmp2589[1], tmp2589[2], tmp2589[3], tmp2589[4], tmp2589[5], tmp2589[6], tmp2589[7]};
    assign tmp1956 = {tmp1955[0], tmp1955[1], tmp1955[2], tmp1955[3], tmp1955[4], tmp1955[5], tmp1955[6], tmp1955[7]};
    assign tmp1561 = {tmp1560, tmp1500};
    assign tmp2399 = tmp2470;
    assign tmp356 = tmp515;
        assign tmp171 = mem_1[b4_w27];
    assign tmp1686 = tmp1682 ^ tmp1685;
        assign tmp2065 = mem_1[tmp2033];
    assign tmp2854 = tmp2850 ^ tmp2853;
    assign tmp394 = tmp390 ^ tmp393;
        assign tmp2704 = mem_3[tmp2672];
        assign tmp1091 = mem_4[tmp927];
    assign tmp2201 = {tmp2200[0], tmp2200[1], tmp2200[2], tmp2200[3], tmp2200[4], tmp2200[5], tmp2200[6], tmp2200[7]};
    assign tmp490 = tmp486 ^ tmp489;
        assign tmp600 = mem_1[tmp568];
    assign c1_w3 = tmp18;
    assign tmp2600 = {tmp2599, tmp2393};
    assign input_wire_10 = temp_35;
        assign tmp1760 = mem_1[tmp1728];
    assign tmp969 = {tmp968[0], tmp968[1], tmp968[2], tmp968[3], tmp968[4], tmp968[5], tmp968[6], tmp968[7]};
    assign tmp538 = tmp534 ^ tmp537;
    assign tmp1331 = {const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0, const1330_0};
    assign c2_w3 = tmp19;
        assign tmp433 = mem_4[tmp335];
    assign tmp1142 = {temp_12[112], temp_12[113], temp_12[114], temp_12[115], temp_12[116], temp_12[117], temp_12[118], temp_12[119]};
    assign tmp2218 = {const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0, const2217_0};
    assign tmp1538 = tmp1534 ^ tmp1537;
    assign temp_13 = tmp1189;
        assign tmp1186 = mem_1[tmp1154];
    assign tmp348 = tmp419;
    assign a1_w15 = tmp84;
    assign tmp163 = {a2_w27, a3_w27, a4_w27, a1_w27};
    assign tmp2685 = {temp_34[16], temp_34[17], temp_34[18], temp_34[19], temp_34[20], temp_34[21], temp_34[22], temp_34[23]};
    assign tmp869 = tmp885;
    assign tmp637 = tmp664;
    assign tmp760 = {tmp759[0], tmp759[1], tmp759[2], tmp759[3], tmp759[4], tmp759[5], tmp759[6], tmp759[7]};
    assign rc3_w3 = const26_0;
        assign tmp589 = mem_1[tmp557];
    assign tmp2629 = tmp2645;
    assign tmp67 = {shifted_w11[0], shifted_w11[1], shifted_w11[2], shifted_w11[3], shifted_w11[4], shifted_w11[5], shifted_w11[6], shifted_w11[7]};
    assign rc2_w35 = const225_0;
    assign tmp1787 = {temp_21[32], temp_21[33], temp_21[34], temp_21[35], temp_21[36], temp_21[37], temp_21[38], temp_21[39]};
        assign tmp93 = mem_1[b1_w15];
    assign tmp2091 = {temp_26[80], temp_26[81], temp_26[82], temp_26[83], temp_26[84], temp_26[85], temp_26[86], temp_26[87]};
    assign tmp2461 = tmp2459 ^ tmp2460;
        assign tmp2067 = mem_1[tmp2035];
    assign tmp1337 = tmp1335 ^ tmp1336;
    assign tmp628 = {temp_6[64], temp_6[65], temp_6[66], temp_6[67], temp_6[68], temp_6[69], temp_6[70], temp_6[71]};
    assign c3_w7 = tmp45;
    assign tmp2864 = {const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0, const2863_0};
    assign tmp522 = tmp518 ^ tmp521;
        assign tmp1311 = mem_3[tmp1213];
    assign tmp2739 = {tmp2738[0], tmp2738[1], tmp2738[2], tmp2738[3], tmp2738[4], tmp2738[5], tmp2738[6], tmp2738[7]};
    assign tmp337 = {temp_2[48], temp_2[49], temp_2[50], temp_2[51], temp_2[52], temp_2[53], temp_2[54], temp_2[55]};
    assign tmp236 = {tmp233[8], tmp233[9], tmp233[10], tmp233[11], tmp233[12], tmp233[13], tmp233[14], tmp233[15]};
        assign tmp665 = mem_3[tmp622];
    assign tmp1576 = {const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0, const1575_0};
    assign tmp2049 = tmp2065;
    assign tmp853 = {temp_8[80], temp_8[81], temp_8[82], temp_8[83], temp_8[84], temp_8[85], temp_8[86], temp_8[87]};
    assign temp_5 = tmp603;
    assign tmp2897 = {expanded_key[128], expanded_key[129], expanded_key[130], expanded_key[131], expanded_key[132], expanded_key[133], expanded_key[134], expanded_key[135], expanded_key[136], expanded_key[137], expanded_key[138], expanded_key[139], expanded_key[140], expanded_key[141], expanded_key[142], expanded_key[143], expanded_key[144], expanded_key[145], expanded_key[146], expanded_key[147], expanded_key[148], expanded_key[149], expanded_key[150], expanded_key[151], expanded_key[152], expanded_key[153], expanded_key[154], expanded_key[155], expanded_key[156], expanded_key[157], expanded_key[158], expanded_key[159], expanded_key[160], expanded_key[161], expanded_key[162], expanded_key[163], expanded_key[164], expanded_key[165], expanded_key[166], expanded_key[167], expanded_key[168], expanded_key[169], expanded_key[170], expanded_key[171], expanded_key[172], expanded_key[173], expanded_key[174], expanded_key[175], expanded_key[176], expanded_key[177], expanded_key[178], expanded_key[179], expanded_key[180], expanded_key[181], expanded_key[182], expanded_key[183], expanded_key[184], expanded_key[185], expanded_key[186], expanded_key[187], expanded_key[188], expanded_key[189], expanded_key[190], expanded_key[191], expanded_key[192], expanded_key[193], expanded_key[194], expanded_key[195], expanded_key[196], expanded_key[197], expanded_key[198], expanded_key[199], expanded_key[200], expanded_key[201], expanded_key[202], expanded_key[203], expanded_key[204], expanded_key[205], expanded_key[206], expanded_key[207], expanded_key[208], expanded_key[209], expanded_key[210], expanded_key[211], expanded_key[212], expanded_key[213], expanded_key[214], expanded_key[215], expanded_key[216], expanded_key[217], expanded_key[218], expanded_key[219], expanded_key[220], expanded_key[221], expanded_key[222], expanded_key[223], expanded_key[224], expanded_key[225], expanded_key[226], expanded_key[227], expanded_key[228], expanded_key[229], expanded_key[230], expanded_key[231], expanded_key[232], expanded_key[233], expanded_key[234], expanded_key[235], expanded_key[236], expanded_key[237], expanded_key[238], expanded_key[239], expanded_key[240], expanded_key[241], expanded_key[242], expanded_key[243], expanded_key[244], expanded_key[245], expanded_key[246], expanded_key[247], expanded_key[248], expanded_key[249], expanded_key[250], expanded_key[251], expanded_key[252], expanded_key[253], expanded_key[254], expanded_key[255]};
    assign tmp122 = {c1_w19, c2_w19, c3_w19, c4_w19};
    assign tmp871 = tmp887;
    assign tmp525 = {tmp524, tmp340};
    assign tmp1137 = {tmp1136[0], tmp1136[1], tmp1136[2], tmp1136[3], tmp1136[4], tmp1136[5], tmp1136[6], tmp1136[7]};
        assign tmp96 = mem_1[b4_w15];
    assign tmp799 = tmp797 ^ tmp798;
    assign tmp2846 = tmp2842 ^ tmp2845;
    assign tmp2152 = tmp2148 ^ tmp2151;
    assign tmp2501 = tmp2497 ^ tmp2500;
    assign tmp113 = {a2_w19, a3_w19, a4_w19, a1_w19};
    assign tmp1209 = {temp_14[104], temp_14[105], temp_14[106], temp_14[107], temp_14[108], temp_14[109], temp_14[110], temp_14[111]};
    assign tmp1738 = {temp_20[32], temp_20[33], temp_20[34], temp_20[35], temp_20[36], temp_20[37], temp_20[38], temp_20[39]};
    assign tmp2177 = {tmp2176[0], tmp2176[1], tmp2176[2], tmp2176[3], tmp2176[4], tmp2176[5], tmp2176[6], tmp2176[7]};
    assign tmp1208 = {temp_14[112], temp_14[113], temp_14[114], temp_14[115], temp_14[116], temp_14[117], temp_14[118], temp_14[119]};
    assign tmp1822 = tmp1992;
    assign tmp2913 = {temp_36[8], temp_36[9], temp_36[10], temp_36[11], temp_36[12], temp_36[13], temp_36[14], temp_36[15]};
    assign tmp1160 = tmp1176;
    assign tmp238 = {a2_w39, a3_w39, a4_w39, a1_w39};
    assign tmp1222 = {temp_14[0], temp_14[1], temp_14[2], temp_14[3], temp_14[4], temp_14[5], temp_14[6], temp_14[7]};
    assign tmp2917 = tmp2933;
    assign tmp2467 = {const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0, const2466_0};
    assign tmp1698 = tmp1694 ^ tmp1697;
        assign tmp2053 = mem_1[tmp2021];
    assign xor_w39 = tmp254;
    assign tmp2727 = {tmp2726[0], tmp2726[1], tmp2726[2], tmp2726[3], tmp2726[4], tmp2726[5], tmp2726[6], tmp2726[7]};
        assign tmp654 = mem_4[tmp622];
    assign tmp1911 = tmp1909 ^ tmp1910;
    assign tmp1961 = {const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0, const1960_0};
    assign w5 = tmp31;
    assign tmp2171 = {tmp2170, tmp2092};
    assign tmp1937 = {const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0, const1936_0};
    assign tmp2720 = {const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0, const2719_0};
    assign c3_w39 = tmp245;
    assign tmp2126 = {const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0, const2125_0};
    assign tmp2374 = {temp_29[24], temp_29[25], temp_29[26], temp_29[27], temp_29[28], temp_29[29], temp_29[30], temp_29[31]};
    assign b2_w31 = tmp190;
    assign tmp2400 = tmp2482;
    assign tmp573 = tmp589;
    assign tmp1932 = {tmp1931[0], tmp1931[1], tmp1931[2], tmp1931[3], tmp1931[4], tmp1931[5], tmp1931[6], tmp1931[7]};
    assign xor_w23 = tmp154;
    assign tmp1010 = {const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0, const1009_0};
    assign rc2_w3 = const25_0;
        assign tmp1981 = mem_3[tmp1806];
    assign tmp1082 = {const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0, const1081_0};
    assign tmp1124 = tmp1120 ^ tmp1123;
    assign c4_w23 = tmp146;
    assign tmp707 = tmp703 ^ tmp706;
    assign tmp34 = {w7[24], w7[25], w7[26], w7[27], w7[28], w7[29], w7[30], w7[31]};
    assign tmp31 = w4 ^ w1;
    assign tmp1444 = {temp_16[40], temp_16[41], temp_16[42], temp_16[43], temp_16[44], temp_16[45], temp_16[46], temp_16[47]};
    assign tmp1257 = tmp1253 ^ tmp1256;
        assign tmp1187 = mem_1[tmp1155];
        assign tmp2130 = mem_3[tmp2087];
    assign tmp395 = {tmp394[0], tmp394[1], tmp394[2], tmp394[3], tmp394[4], tmp394[5], tmp394[6], tmp394[7]};
    assign tmp1272 = {tmp1271, tmp1208};
    assign tmp916 = {temp_10[104], temp_10[105], temp_10[106], temp_10[107], temp_10[108], temp_10[109], temp_10[110], temp_10[111]};
    assign tmp2243 = {tmp2242, tmp2094};
        assign tmp1478 = mem_1[tmp1446];
        assign tmp99 = mem_2[const98_4];
        assign tmp890 = mem_1[tmp858];
    assign tmp1855 = tmp1851 ^ tmp1854;
    assign tmp2630 = tmp2646;
    assign tmp2320 = {temp_28[64], temp_28[65], temp_28[66], temp_28[67], temp_28[68], temp_28[69], temp_28[70], temp_28[71]};
    assign tmp2103 = tmp2141;
    assign tmp2500 = {tmp2499, tmp2384};
    assign tmp2903 = {temp_36[88], temp_36[89], temp_36[90], temp_36[91], temp_36[92], temp_36[93], temp_36[94], temp_36[95]};
    assign tmp1519 = tmp1579;
    assign tmp405 = {tmp404, tmp330};
    assign tmp1509 = {temp_18[48], temp_18[49], temp_18[50], temp_18[51], temp_18[52], temp_18[53], temp_18[54], temp_18[55]};
    assign tmp1851 = tmp1849 ^ tmp1850;
    assign tmp2911 = {temp_36[24], temp_36[25], temp_36[26], temp_36[27], temp_36[28], temp_36[29], temp_36[30], temp_36[31]};
    assign tmp2504 = {tmp2503, tmp2385};
    assign tmp1432 = {expanded_key[768], expanded_key[769], expanded_key[770], expanded_key[771], expanded_key[772], expanded_key[773], expanded_key[774], expanded_key[775], expanded_key[776], expanded_key[777], expanded_key[778], expanded_key[779], expanded_key[780], expanded_key[781], expanded_key[782], expanded_key[783], expanded_key[784], expanded_key[785], expanded_key[786], expanded_key[787], expanded_key[788], expanded_key[789], expanded_key[790], expanded_key[791], expanded_key[792], expanded_key[793], expanded_key[794], expanded_key[795], expanded_key[796], expanded_key[797], expanded_key[798], expanded_key[799], expanded_key[800], expanded_key[801], expanded_key[802], expanded_key[803], expanded_key[804], expanded_key[805], expanded_key[806], expanded_key[807], expanded_key[808], expanded_key[809], expanded_key[810], expanded_key[811], expanded_key[812], expanded_key[813], expanded_key[814], expanded_key[815], expanded_key[816], expanded_key[817], expanded_key[818], expanded_key[819], expanded_key[820], expanded_key[821], expanded_key[822], expanded_key[823], expanded_key[824], expanded_key[825], expanded_key[826], expanded_key[827], expanded_key[828], expanded_key[829], expanded_key[830], expanded_key[831], expanded_key[832], expanded_key[833], expanded_key[834], expanded_key[835], expanded_key[836], expanded_key[837], expanded_key[838], expanded_key[839], expanded_key[840], expanded_key[841], expanded_key[842], expanded_key[843], expanded_key[844], expanded_key[845], expanded_key[846], expanded_key[847], expanded_key[848], expanded_key[849], expanded_key[850], expanded_key[851], expanded_key[852], expanded_key[853], expanded_key[854], expanded_key[855], expanded_key[856], expanded_key[857], expanded_key[858], expanded_key[859], expanded_key[860], expanded_key[861], expanded_key[862], expanded_key[863], expanded_key[864], expanded_key[865], expanded_key[866], expanded_key[867], expanded_key[868], expanded_key[869], expanded_key[870], expanded_key[871], expanded_key[872], expanded_key[873], expanded_key[874], expanded_key[875], expanded_key[876], expanded_key[877], expanded_key[878], expanded_key[879], expanded_key[880], expanded_key[881], expanded_key[882], expanded_key[883], expanded_key[884], expanded_key[885], expanded_key[886], expanded_key[887], expanded_key[888], expanded_key[889], expanded_key[890], expanded_key[891], expanded_key[892], expanded_key[893], expanded_key[894], expanded_key[895]};
    assign tmp1139 = {expanded_key[896], expanded_key[897], expanded_key[898], expanded_key[899], expanded_key[900], expanded_key[901], expanded_key[902], expanded_key[903], expanded_key[904], expanded_key[905], expanded_key[906], expanded_key[907], expanded_key[908], expanded_key[909], expanded_key[910], expanded_key[911], expanded_key[912], expanded_key[913], expanded_key[914], expanded_key[915], expanded_key[916], expanded_key[917], expanded_key[918], expanded_key[919], expanded_key[920], expanded_key[921], expanded_key[922], expanded_key[923], expanded_key[924], expanded_key[925], expanded_key[926], expanded_key[927], expanded_key[928], expanded_key[929], expanded_key[930], expanded_key[931], expanded_key[932], expanded_key[933], expanded_key[934], expanded_key[935], expanded_key[936], expanded_key[937], expanded_key[938], expanded_key[939], expanded_key[940], expanded_key[941], expanded_key[942], expanded_key[943], expanded_key[944], expanded_key[945], expanded_key[946], expanded_key[947], expanded_key[948], expanded_key[949], expanded_key[950], expanded_key[951], expanded_key[952], expanded_key[953], expanded_key[954], expanded_key[955], expanded_key[956], expanded_key[957], expanded_key[958], expanded_key[959], expanded_key[960], expanded_key[961], expanded_key[962], expanded_key[963], expanded_key[964], expanded_key[965], expanded_key[966], expanded_key[967], expanded_key[968], expanded_key[969], expanded_key[970], expanded_key[971], expanded_key[972], expanded_key[973], expanded_key[974], expanded_key[975], expanded_key[976], expanded_key[977], expanded_key[978], expanded_key[979], expanded_key[980], expanded_key[981], expanded_key[982], expanded_key[983], expanded_key[984], expanded_key[985], expanded_key[986], expanded_key[987], expanded_key[988], expanded_key[989], expanded_key[990], expanded_key[991], expanded_key[992], expanded_key[993], expanded_key[994], expanded_key[995], expanded_key[996], expanded_key[997], expanded_key[998], expanded_key[999], expanded_key[1000], expanded_key[1001], expanded_key[1002], expanded_key[1003], expanded_key[1004], expanded_key[1005], expanded_key[1006], expanded_key[1007], expanded_key[1008], expanded_key[1009], expanded_key[1010], expanded_key[1011], expanded_key[1012], expanded_key[1013], expanded_key[1014], expanded_key[1015], expanded_key[1016], expanded_key[1017], expanded_key[1018], expanded_key[1019], expanded_key[1020], expanded_key[1021], expanded_key[1022], expanded_key[1023]};
    assign tmp751 = tmp749 ^ tmp750;
    assign tmp996 = tmp994 ^ tmp995;
    assign tmp371 = {tmp370[0], tmp370[1], tmp370[2], tmp370[3], tmp370[4], tmp370[5], tmp370[6], tmp370[7]};
    assign tmp1574 = tmp1570 ^ tmp1573;
    assign tmp286 = tmp302;
        assign tmp2824 = mem_3[tmp2682];
    assign tmp2234 = {const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0, const2233_0};
    assign tmp2025 = {temp_24[80], temp_24[81], temp_24[82], temp_24[83], temp_24[84], temp_24[85], temp_24[86], temp_24[87]};
        assign tmp143 = mem_1[b1_w23];
        assign tmp2299 = mem_4[tmp2098];
    assign tmp1918 = {tmp1917, tmp1799};
    assign tmp2377 = {temp_29[0], temp_29[1], temp_29[2], temp_29[3], temp_29[4], temp_29[5], temp_29[6], temp_29[7]};
    assign tmp129 = concat_w19 ^ substituted_w19;
    assign tmp2547 = {const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0, const2546_0};
    assign tmp1591 = {tmp1590[0], tmp1590[1], tmp1590[2], tmp1590[3], tmp1590[4], tmp1590[5], tmp1590[6], tmp1590[7]};
    assign tmp1512 = {temp_18[24], temp_18[25], temp_18[26], temp_18[27], temp_18[28], temp_18[29], temp_18[30], temp_18[31]};
    assign tmp332 = {temp_2[88], temp_2[89], temp_2[90], temp_2[91], temp_2[92], temp_2[93], temp_2[94], temp_2[95]};
    assign tmp1207 = {temp_14[120], temp_14[121], temp_14[122], temp_14[123], temp_14[124], temp_14[125], temp_14[126], temp_14[127]};
    assign tmp1229 = tmp1322;
        assign tmp444 = mem_3[tmp335];
    assign tmp78 = {rc1_w11, rc2_w11, rc3_w11, rc4_w11};
    assign tmp2965 = {expanded_key[0], expanded_key[1], expanded_key[2], expanded_key[3], expanded_key[4], expanded_key[5], expanded_key[6], expanded_key[7], expanded_key[8], expanded_key[9], expanded_key[10], expanded_key[11], expanded_key[12], expanded_key[13], expanded_key[14], expanded_key[15], expanded_key[16], expanded_key[17], expanded_key[18], expanded_key[19], expanded_key[20], expanded_key[21], expanded_key[22], expanded_key[23], expanded_key[24], expanded_key[25], expanded_key[26], expanded_key[27], expanded_key[28], expanded_key[29], expanded_key[30], expanded_key[31], expanded_key[32], expanded_key[33], expanded_key[34], expanded_key[35], expanded_key[36], expanded_key[37], expanded_key[38], expanded_key[39], expanded_key[40], expanded_key[41], expanded_key[42], expanded_key[43], expanded_key[44], expanded_key[45], expanded_key[46], expanded_key[47], expanded_key[48], expanded_key[49], expanded_key[50], expanded_key[51], expanded_key[52], expanded_key[53], expanded_key[54], expanded_key[55], expanded_key[56], expanded_key[57], expanded_key[58], expanded_key[59], expanded_key[60], expanded_key[61], expanded_key[62], expanded_key[63], expanded_key[64], expanded_key[65], expanded_key[66], expanded_key[67], expanded_key[68], expanded_key[69], expanded_key[70], expanded_key[71], expanded_key[72], expanded_key[73], expanded_key[74], expanded_key[75], expanded_key[76], expanded_key[77], expanded_key[78], expanded_key[79], expanded_key[80], expanded_key[81], expanded_key[82], expanded_key[83], expanded_key[84], expanded_key[85], expanded_key[86], expanded_key[87], expanded_key[88], expanded_key[89], expanded_key[90], expanded_key[91], expanded_key[92], expanded_key[93], expanded_key[94], expanded_key[95], expanded_key[96], expanded_key[97], expanded_key[98], expanded_key[99], expanded_key[100], expanded_key[101], expanded_key[102], expanded_key[103], expanded_key[104], expanded_key[105], expanded_key[106], expanded_key[107], expanded_key[108], expanded_key[109], expanded_key[110], expanded_key[111], expanded_key[112], expanded_key[113], expanded_key[114], expanded_key[115], expanded_key[116], expanded_key[117], expanded_key[118], expanded_key[119], expanded_key[120], expanded_key[121], expanded_key[122], expanded_key[123], expanded_key[124], expanded_key[125], expanded_key[126], expanded_key[127]};
    assign tmp498 = tmp494 ^ tmp497;
    assign tmp343 = {temp_2[0], temp_2[1], temp_2[2], temp_2[3], temp_2[4], temp_2[5], temp_2[6], temp_2[7]};
    assign tmp110 = {tmp108[16], tmp108[17], tmp108[18], tmp108[19], tmp108[20], tmp108[21], tmp108[22], tmp108[23]};
        assign tmp2203 = mem_4[tmp2090];
    assign tmp2086 = {temp_26[120], temp_26[121], temp_26[122], temp_26[123], temp_26[124], temp_26[125], temp_26[126], temp_26[127]};
    assign tmp1754 = tmp1770;
    assign tmp2010 = {tmp2009, tmp1806};
    assign tmp1989 = {const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0, const1988_0};
    assign tmp500 = {const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0, const499_0};
        assign tmp2471 = mem_3[tmp2384];
        assign tmp1772 = mem_1[tmp1740];
        assign tmp2251 = mem_4[tmp2094];
    assign tmp272 = {new_state[40], new_state[41], new_state[42], new_state[43], new_state[44], new_state[45], new_state[46], new_state[47]};
    assign tmp1550 = tmp1546 ^ tmp1549;
    assign tmp621 = {temp_6[120], temp_6[121], temp_6[122], temp_6[123], temp_6[124], temp_6[125], temp_6[126], temp_6[127]};
    assign tmp616 = {temp_5[24], temp_5[25], temp_5[26], temp_5[27], temp_5[28], temp_5[29], temp_5[30], temp_5[31]};
    assign c1_w27 = tmp168;
    assign tmp1192 = {temp_13[104], temp_13[105], temp_13[106], temp_13[107], temp_13[108], temp_13[109], temp_13[110], temp_13[111]};
    assign tmp1820 = tmp1968;
    assign tmp2871 = {tmp2870[0], tmp2870[1], tmp2870[2], tmp2870[3], tmp2870[4], tmp2870[5], tmp2870[6], tmp2870[7]};
        assign tmp1251 = mem_3[tmp1208];
    assign tmp1154 = {temp_12[16], temp_12[17], temp_12[18], temp_12[19], temp_12[20], temp_12[21], temp_12[22], temp_12[23]};
    assign tmp2695 = tmp2799;
    assign rc1_w39 = tmp249;
    assign tmp1742 = {temp_20[0], temp_20[1], temp_20[2], temp_20[3], temp_20[4], temp_20[5], temp_20[6], temp_20[7]};
    assign tmp2497 = tmp2495 ^ tmp2496;
    assign tmp2811 = {tmp2810[0], tmp2810[1], tmp2810[2], tmp2810[3], tmp2810[4], tmp2810[5], tmp2810[6], tmp2810[7]};
    assign tmp183 = tmp182 ^ tmp158;
    assign tmp489 = {tmp488, tmp337};
    assign tmp1791 = {temp_21[0], temp_21[1], temp_21[2], temp_21[3], temp_21[4], temp_21[5], temp_21[6], temp_21[7]};
    assign tmp1991 = tmp1987 ^ tmp1990;
    assign tmp1219 = {temp_14[24], temp_14[25], temp_14[26], temp_14[27], temp_14[28], temp_14[29], temp_14[30], temp_14[31]};
    assign a1_w23 = tmp134;
        assign tmp797 = mem_3[tmp633];
    assign tmp622 = {temp_6[112], temp_6[113], temp_6[114], temp_6[115], temp_6[116], temp_6[117], temp_6[118], temp_6[119]};
    assign tmp1881 = {const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0, const1880_0};
    assign tmp577 = tmp593;
    assign tmp1627 = {tmp1626[0], tmp1626[1], tmp1626[2], tmp1626[3], tmp1626[4], tmp1626[5], tmp1626[6], tmp1626[7]};
    assign tmp1585 = {tmp1584, tmp1506};
    assign tmp2655 = {temp_33[120], temp_33[121], temp_33[122], temp_33[123], temp_33[124], temp_33[125], temp_33[126], temp_33[127]};
    assign tmp1853 = {const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0, const1852_0};
    assign tmp944 = tmp1125;
    assign tmp1644 = {const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0, const1643_0};
    assign tmp2402 = tmp2506;
        assign tmp2214 = mem_3[tmp2094];
    assign tmp1905 = {const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0, const1904_0};
    assign tmp474 = tmp470 ^ tmp473;
    assign tmp2899 = {temp_36[120], temp_36[121], temp_36[122], temp_36[123], temp_36[124], temp_36[125], temp_36[126], temp_36[127]};
    assign tmp1201 = {temp_13[32], temp_13[33], temp_13[34], temp_13[35], temp_13[36], temp_13[37], temp_13[38], temp_13[39]};
    assign tmp1810 = tmp1848;
    assign tmp446 = tmp444 ^ tmp445;
    assign tmp1962 = {tmp1961, tmp1802};
    assign tmp2926 = tmp2942;
    assign tmp2573 = tmp2569 ^ tmp2572;
    assign tmp2115 = tmp2285;
    assign tmp1346 = {tmp1345[0], tmp1345[1], tmp1345[2], tmp1345[3], tmp1345[4], tmp1345[5], tmp1345[6], tmp1345[7]};
    assign tmp964 = tmp960 ^ tmp963;
    assign tmp1753 = tmp1769;
    assign tmp950 = {const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0, const949_0};
    assign tmp877 = tmp893;
    assign tmp1925 = {const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0, const1924_0};
    assign tmp1613 = {tmp1612, tmp1505};
    assign tmp838 = {tmp837, tmp634};
    assign tmp986 = {const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0, const985_0};
    assign tmp1668 = {const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0, const1667_0};
    assign tmp554 = temp_3 ^ tmp553;
    assign tmp2294 = {const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0, const2293_0};
    assign tmp191 = {shifted_w31[8], shifted_w31[9], shifted_w31[10], shifted_w31[11], shifted_w31[12], shifted_w31[13], shifted_w31[14], shifted_w31[15]};
        assign tmp1175 = mem_1[tmp1143];
    assign tmp1517 = tmp1555;
    assign tmp1112 = tmp1108 ^ tmp1111;
    assign tmp2516 = {tmp2515, tmp2390};
        assign tmp2942 = mem_1[tmp2910];
    assign tmp2823 = {tmp2822[0], tmp2822[1], tmp2822[2], tmp2822[3], tmp2822[4], tmp2822[5], tmp2822[6], tmp2822[7]};
    assign tmp917 = {temp_10[96], temp_10[97], temp_10[98], temp_10[99], temp_10[100], temp_10[101], temp_10[102], temp_10[103]};
    assign tmp1143 = {temp_12[104], temp_12[105], temp_12[106], temp_12[107], temp_12[108], temp_12[109], temp_12[110], temp_12[111]};
    assign tmp1092 = tmp1090 ^ tmp1091;
    assign tmp1050 = {const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0, const1049_0};
    assign tmp935 = tmp1017;
    assign tmp2605 = temp_31 ^ tmp2604;
    assign tmp911 = {temp_9[8], temp_9[9], temp_9[10], temp_9[11], temp_9[12], temp_9[13], temp_9[14], temp_9[15]};
    assign tmp2915 = tmp2931;
    assign tmp1860 = {tmp1859[0], tmp1859[1], tmp1859[2], tmp1859[3], tmp1859[4], tmp1859[5], tmp1859[6], tmp1859[7]};
    assign tmp2326 = {temp_28[16], temp_28[17], temp_28[18], temp_28[19], temp_28[20], temp_28[21], temp_28[22], temp_28[23]};
    assign tmp2188 = tmp2184 ^ tmp2187;
        assign tmp1958 = mem_4[tmp1801];
    assign tmp1739 = {temp_20[24], temp_20[25], temp_20[26], temp_20[27], temp_20[28], temp_20[29], temp_20[30], temp_20[31]};
    assign tmp1329 = tmp1325 ^ tmp1328;
    assign tmp312 = {temp_1[112], temp_1[113], temp_1[114], temp_1[115], temp_1[116], temp_1[117], temp_1[118], temp_1[119]};
        assign tmp2932 = mem_1[tmp2900];
        assign tmp1185 = mem_1[tmp1153];
        assign tmp2765 = mem_4[tmp2678];
    assign tmp2676 = {temp_34[88], temp_34[89], temp_34[90], temp_34[91], temp_34[92], temp_34[93], temp_34[94], temp_34[95]};
    assign tmp230 = tmp205 ^ xor_w35;
    assign tmp2596 = {tmp2595, tmp2392};
        assign tmp1475 = mem_1[tmp1443];
    assign tmp350 = tmp443;
    assign tmp2806 = tmp2802 ^ tmp2805;
    assign tmp107 = tmp106 ^ tmp82;
    assign tmp2200 = tmp2196 ^ tmp2199;
    assign tmp2540 = {tmp2539, tmp2388};
    assign tmp706 = {tmp705, tmp627};
    assign tmp930 = tmp957;
    assign tmp2022 = {temp_24[104], temp_24[105], temp_24[106], temp_24[107], temp_24[108], temp_24[109], temp_24[110], temp_24[111]};
    assign tmp711 = tmp707 ^ tmp710;
        assign tmp1323 = mem_3[tmp1214];
        assign tmp196 = mem_1[b4_w31];
        assign tmp822 = mem_4[tmp636];
    assign tmp2403 = tmp2518;
        assign tmp516 = mem_3[tmp341];
    assign tmp1489 = {temp_17[72], temp_17[73], temp_17[74], temp_17[75], temp_17[76], temp_17[77], temp_17[78], temp_17[79]};
    assign tmp319 = {temp_1[56], temp_1[57], temp_1[58], temp_1[59], temp_1[60], temp_1[61], temp_1[62], temp_1[63]};
    assign tmp2453 = tmp2449 ^ tmp2452;
    assign tmp87 = {tmp83[0], tmp83[1], tmp83[2], tmp83[3], tmp83[4], tmp83[5], tmp83[6], tmp83[7]};
    assign tmp32 = w5 ^ w2;
        assign tmp2459 = mem_3[tmp2383];
    assign tmp2909 = {temp_36[40], temp_36[41], temp_36[42], temp_36[43], temp_36[44], temp_36[45], temp_36[46], temp_36[47]};
    assign tmp2742 = tmp2740 ^ tmp2741;
    assign tmp790 = {tmp789, tmp630};
    assign tmp1053 = {tmp1052[0], tmp1052[1], tmp1052[2], tmp1052[3], tmp1052[4], tmp1052[5], tmp1052[6], tmp1052[7]};
    assign tmp2421 = tmp2417 ^ tmp2420;
    assign tmp1642 = tmp1640 ^ tmp1641;
    assign tmp1385 = tmp1383 ^ tmp1384;
        assign tmp1347 = mem_3[tmp1216];
    assign tmp1077 = {tmp1076[0], tmp1076[1], tmp1076[2], tmp1076[3], tmp1076[4], tmp1076[5], tmp1076[6], tmp1076[7]};
    assign tmp2208 = tmp2204 ^ tmp2207;
    assign tmp922 = {temp_10[56], temp_10[57], temp_10[58], temp_10[59], temp_10[60], temp_10[61], temp_10[62], temp_10[63]};
        assign tmp1288 = mem_4[tmp1212];
    assign tmp508 = {const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0, const507_0};
    assign tmp2220 = tmp2216 ^ tmp2219;
    assign shifted_w27 = tmp163;
        assign tmp1276 = mem_4[tmp1207];
    assign tmp2081 = {temp_25[24], temp_25[25], temp_25[26], temp_25[27], temp_25[28], temp_25[29], temp_25[30], temp_25[31]};
    assign tmp1799 = {temp_22[72], temp_22[73], temp_22[74], temp_22[75], temp_22[76], temp_22[77], temp_22[78], temp_22[79]};
    assign a4_w15 = tmp87;
    assign tmp820 = {tmp819[0], tmp819[1], tmp819[2], tmp819[3], tmp819[4], tmp819[5], tmp819[6], tmp819[7]};
    assign tmp188 = {a2_w31, a3_w31, a4_w31, a1_w31};
        assign tmp2063 = mem_1[tmp2031];
    assign b3_w27 = tmp166;
        assign tmp1018 = mem_3[tmp920];
    assign tmp2798 = tmp2794 ^ tmp2797;
    assign tmp1376 = {tmp1375, tmp1216};
    assign tmp2134 = {const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0, const2133_0};
    assign tmp1931 = tmp1927 ^ tmp1930;
    assign tmp207 = tmp206 ^ tmp182;
    assign tmp700 = {tmp699[0], tmp699[1], tmp699[2], tmp699[3], tmp699[4], tmp699[5], tmp699[6], tmp699[7]};
        assign tmp2873 = mem_4[tmp2687];
    assign tmp1411 = {const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0, const1410_0};
    assign tmp687 = tmp683 ^ tmp686;
        assign tmp983 = mem_4[tmp914];
    assign substituted_w19 = tmp122;
        assign tmp2741 = mem_4[tmp2672];
    assign tmp166 = {shifted_w27[8], shifted_w27[9], shifted_w27[10], shifted_w27[11], shifted_w27[12], shifted_w27[13], shifted_w27[14], shifted_w27[15]};
    assign tmp1598 = tmp1594 ^ tmp1597;
    assign tmp1803 = {temp_22[40], temp_22[41], temp_22[42], temp_22[43], temp_22[44], temp_22[45], temp_22[46], temp_22[47]};
    assign tmp962 = {const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0, const961_0};
        assign tmp70 = mem_1[b3_w11];
    assign tmp1674 = tmp1670 ^ tmp1673;
    assign tmp2248 = tmp2244 ^ tmp2247;
    assign tmp82 = tmp81 ^ tmp57;
    assign tmp641 = tmp712;
    assign tmp1373 = tmp1371 ^ tmp1372;
    assign tmp2624 = tmp2640;
    assign xor_w31 = tmp204;
    assign tmp2696 = tmp2811;
    assign tmp1212 = {temp_14[80], temp_14[81], temp_14[82], temp_14[83], temp_14[84], temp_14[85], temp_14[86], temp_14[87]};
    assign tmp1450 = tmp1466;
        assign tmp244 = mem_1[b2_w39];
        assign tmp2729 = mem_4[tmp2675];
    assign tmp1777 = {temp_21[112], temp_21[113], temp_21[114], temp_21[115], temp_21[116], temp_21[117], temp_21[118], temp_21[119]};
    assign tmp2102 = tmp2129;
        assign tmp2066 = mem_1[tmp2034];
    assign tmp2689 = tmp2727;
    assign tmp284 = tmp300;
    assign tmp555 = {temp_4[120], temp_4[121], temp_4[122], temp_4[123], temp_4[124], temp_4[125], temp_4[126], temp_4[127]};
    assign tmp261 = aes_plaintext ^ tmp260;
    assign tmp401 = {tmp400, tmp329};
    assign tmp1758 = tmp1774;
    assign tmp1391 = {const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0, const1390_0};
        assign tmp702 = mem_4[tmp626];
    assign tmp1083 = {tmp1082, tmp923};
    assign tmp2192 = tmp2190 ^ tmp2191;
    assign tmp2822 = tmp2818 ^ tmp2821;
    assign tmp1908 = {tmp1907[0], tmp1907[1], tmp1907[2], tmp1907[3], tmp1907[4], tmp1907[5], tmp1907[6], tmp1907[7]};
    assign tmp560 = {temp_4[80], temp_4[81], temp_4[82], temp_4[83], temp_4[84], temp_4[85], temp_4[86], temp_4[87]};
    assign tmp2048 = tmp2064;
        assign tmp249 = mem_2[const248_10];
    assign tmp1813 = tmp1884;
    assign tmp929 = {temp_10[0], temp_10[1], temp_10[2], temp_10[3], temp_10[4], temp_10[5], temp_10[6], temp_10[7]};
    assign tmp2690 = tmp2739;
    assign tmp960 = tmp958 ^ tmp959;
    assign tmp2769 = {tmp2768, tmp2679};
    assign new_10 = tmp2898;
        assign tmp300 = mem_1[tmp268];
    assign tmp865 = tmp881;
    assign tmp2530 = {tmp2529[0], tmp2529[1], tmp2529[2], tmp2529[3], tmp2529[4], tmp2529[5], tmp2529[6], tmp2529[7]};
    assign tmp1293 = tmp1289 ^ tmp1292;
    assign tmp228 = {rc1_w35, rc2_w35, rc3_w35, rc4_w35};
    assign tmp352 = tmp467;
    assign tmp536 = {const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0, const535_0};
    assign tmp2382 = {temp_30[96], temp_30[97], temp_30[98], temp_30[99], temp_30[100], temp_30[101], temp_30[102], temp_30[103]};
    assign tmp1899 = tmp1897 ^ tmp1898;
    assign tmp1680 = {const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0, const1679_0};
    assign tmp2782 = tmp2778 ^ tmp2781;
    assign tmp2033 = {temp_24[16], temp_24[17], temp_24[18], temp_24[19], temp_24[20], temp_24[21], temp_24[22], temp_24[23]};
    assign rc1_w15 = tmp99;
    assign tmp2365 = {temp_29[96], temp_29[97], temp_29[98], temp_29[99], temp_29[100], temp_29[101], temp_29[102], temp_29[103]};
    assign tmp1136 = tmp1132 ^ tmp1135;
    assign tmp557 = {temp_4[104], temp_4[105], temp_4[106], temp_4[107], temp_4[108], temp_4[109], temp_4[110], temp_4[111]};
    assign c4_w31 = tmp196;
    assign tmp2893 = {tmp2892, tmp2686};
    assign tmp454 = tmp450 ^ tmp453;
    assign tmp197 = {c1_w31, c2_w31, c3_w31, c4_w31};
    assign c2_w27 = tmp169;
    assign tmp1669 = {tmp1668, tmp1509};
    assign tmp2132 = tmp2130 ^ tmp2131;
    assign tmp1352 = {tmp1351, tmp1218};
    assign tmp1439 = {temp_16[80], temp_16[81], temp_16[82], temp_16[83], temp_16[84], temp_16[85], temp_16[86], temp_16[87]};
        assign tmp2885 = mem_4[tmp2684];
        assign tmp2555 = mem_3[tmp2391];
        assign tmp21 = mem_1[b4_w3];
    assign tmp2963 = {temp_37[0], temp_37[1], temp_37[2], temp_37[3], temp_37[4], temp_37[5], temp_37[6], temp_37[7]};
    assign tmp2158 = {const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0, const2157_0};
        assign tmp298 = mem_1[tmp266];
    assign tmp482 = tmp480 ^ tmp481;
    assign tmp1014 = {const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0, const1013_0};
    assign tmp1281 = tmp1277 ^ tmp1280;
    assign tmp1446 = {temp_16[24], temp_16[25], temp_16[26], temp_16[27], temp_16[28], temp_16[29], temp_16[30], temp_16[31]};
        assign tmp2937 = mem_1[tmp2905];
    assign tmp2952 = {temp_37[88], temp_37[89], temp_37[90], temp_37[91], temp_37[92], temp_37[93], temp_37[94], temp_37[95]};
    assign temp_23 = tmp2017;
    assign tmp2856 = {const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0, const2855_0};
    assign tmp844 = {tmp843[0], tmp843[1], tmp843[2], tmp843[3], tmp843[4], tmp843[5], tmp843[6], tmp843[7]};
    assign b1_w7 = tmp39;
    assign tmp2068 = {tmp2036, tmp2037, tmp2038, tmp2039, tmp2040, tmp2041, tmp2042, tmp2043, tmp2044, tmp2045, tmp2046, tmp2047, tmp2048, tmp2049, tmp2050, tmp2051};
    assign tmp1678 = tmp1676 ^ tmp1677;
    assign tmp212 = {tmp208[0], tmp208[1], tmp208[2], tmp208[3], tmp208[4], tmp208[5], tmp208[6], tmp208[7]};
    assign tmp658 = {tmp657, tmp623};
    assign tmp723 = tmp719 ^ tmp722;
    assign shifted_w35 = tmp213;
    assign c3_w11 = tmp70;
    assign tmp437 = {tmp436, tmp332};
    assign new_8 = tmp2312;
    assign tmp1497 = {temp_17[8], temp_17[9], temp_17[10], temp_17[11], temp_17[12], temp_17[13], temp_17[14], temp_17[15]};
        assign tmp947 = mem_4[tmp915];
    assign tmp2120 = tmp2118 ^ tmp2119;
    assign tmp1286 = {tmp1285[0], tmp1285[1], tmp1285[2], tmp1285[3], tmp1285[4], tmp1285[5], tmp1285[6], tmp1285[7]};
    assign tmp2104 = tmp2153;
        assign tmp1043 = mem_4[tmp923];
    assign tmp2391 = {temp_30[24], temp_30[25], temp_30[26], temp_30[27], temp_30[28], temp_30[29], temp_30[30], temp_30[31]};
    assign tmp465 = {tmp464, tmp339};
        assign tmp2275 = mem_4[tmp2100];
    assign tmp1666 = tmp1664 ^ tmp1665;
    assign tmp746 = {tmp745, tmp627};
    assign a3_w3 = tmp11;
    assign tmp279 = tmp295;
        assign tmp593 = mem_1[tmp561];
    assign tmp876 = tmp892;
    assign tmp2525 = tmp2521 ^ tmp2524;
    assign tmp1151 = {temp_12[40], temp_12[41], temp_12[42], temp_12[43], temp_12[44], temp_12[45], temp_12[46], temp_12[47]};
    assign tmp2264 = tmp2262 ^ tmp2263;
    assign tmp1808 = {temp_22[0], temp_22[1], temp_22[2], temp_22[3], temp_22[4], temp_22[5], temp_22[6], temp_22[7]};
        assign tmp2764 = mem_3[tmp2677];
        assign tmp19 = mem_1[b2_w3];
    assign c1_w15 = tmp93;
        assign tmp2423 = mem_3[tmp2380];
    assign tmp2786 = tmp2782 ^ tmp2785;
    assign tmp237 = {tmp233[0], tmp233[1], tmp233[2], tmp233[3], tmp233[4], tmp233[5], tmp233[6], tmp233[7]};
    assign tmp2895 = {tmp2894[0], tmp2894[1], tmp2894[2], tmp2894[3], tmp2894[4], tmp2894[5], tmp2894[6], tmp2894[7]};
    assign tmp2814 = tmp2812 ^ tmp2813;
        assign tmp1769 = mem_1[tmp1737];
    assign a1_w3 = tmp9;
    assign tmp452 = {const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0, const451_0};
    assign tmp488 = {const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0, const487_0};
    assign tmp568 = {temp_4[16], temp_4[17], temp_4[18], temp_4[19], temp_4[20], temp_4[21], temp_4[22], temp_4[23]};
    assign tmp2097 = {temp_26[32], temp_26[33], temp_26[34], temp_26[35], temp_26[36], temp_26[37], temp_26[38], temp_26[39]};
    assign tmp1167 = tmp1183;
    assign tmp2883 = {tmp2882[0], tmp2882[1], tmp2882[2], tmp2882[3], tmp2882[4], tmp2882[5], tmp2882[6], tmp2882[7]};
        assign tmp1897 = mem_3[tmp1799];
    assign tmp2612 = {temp_32[72], temp_32[73], temp_32[74], temp_32[75], temp_32[76], temp_32[77], temp_32[78], temp_32[79]};
        assign tmp541 = mem_4[tmp340];
    assign tmp1513 = {temp_18[16], temp_18[17], temp_18[18], temp_18[19], temp_18[20], temp_18[21], temp_18[22], temp_18[23]};
    assign tmp1980 = {tmp1979[0], tmp1979[1], tmp1979[2], tmp1979[3], tmp1979[4], tmp1979[5], tmp1979[6], tmp1979[7]};
    assign tmp1745 = tmp1761;
        assign tmp888 = mem_1[tmp856];
    assign tmp902 = {temp_9[80], temp_9[81], temp_9[82], temp_9[83], temp_9[84], temp_9[85], temp_9[86], temp_9[87]};
        assign tmp2345 = mem_1[tmp2313];
    assign tmp2542 = {tmp2541[0], tmp2541[1], tmp2541[2], tmp2541[3], tmp2541[4], tmp2541[5], tmp2541[6], tmp2541[7]};
    assign rc2_w19 = const125_0;
        assign tmp1545 = mem_4[tmp1502];
    assign tmp292 = tmp308;
    assign tmp431 = {tmp430[0], tmp430[1], tmp430[2], tmp430[3], tmp430[4], tmp430[5], tmp430[6], tmp430[7]};
    assign tmp775 = tmp773 ^ tmp774;
    assign tmp2123 = {tmp2122, tmp2088};
    assign tmp84 = {tmp83[24], tmp83[25], tmp83[26], tmp83[27], tmp83[28], tmp83[29], tmp83[30], tmp83[31]};
    assign tmp694 = {tmp693, tmp622};
    assign tmp1779 = {temp_21[96], temp_21[97], temp_21[98], temp_21[99], temp_21[100], temp_21[101], temp_21[102], temp_21[103]};
        assign tmp2005 = mem_3[tmp1808];
        assign tmp1181 = mem_1[tmp1149];
    assign tmp2242 = {const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0, const2241_0};
    assign tmp1802 = {temp_22[48], temp_22[49], temp_22[50], temp_22[51], temp_22[52], temp_22[53], temp_22[54], temp_22[55]};
    assign tmp1926 = {tmp1925, tmp1803};
    assign a1_w27 = tmp159;
    assign tmp537 = {tmp536, tmp341};
    assign tmp281 = tmp297;
    assign tmp1095 = {tmp1094, tmp928};
    assign tmp293 = tmp309;
    assign tmp2339 = tmp2355;
    assign tmp2240 = tmp2238 ^ tmp2239;
        assign tmp701 = mem_3[tmp625];
        assign tmp94 = mem_1[b2_w15];
    assign tmp1038 = {const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0, const1037_0};
    assign tmp675 = tmp671 ^ tmp674;
    assign temp_30 = tmp2378;
    assign tmp549 = {tmp548, tmp342};
    assign tmp2633 = tmp2649;
    assign tmp1499 = {tmp1483, tmp1488, tmp1493, tmp1498, tmp1487, tmp1492, tmp1497, tmp1486, tmp1491, tmp1496, tmp1485, tmp1490, tmp1495, tmp1484, tmp1489, tmp1494};
        assign tmp220 = mem_1[b3_w35];
    assign tmp1570 = tmp1568 ^ tmp1569;
        assign tmp2567 = mem_3[tmp2392];
    assign tmp1427 = {const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0, const1426_0};
    assign tmp1939 = tmp1935 ^ tmp1938;
    assign tmp2364 = {temp_29[104], temp_29[105], temp_29[106], temp_29[107], temp_29[108], temp_29[109], temp_29[110], temp_29[111]};
    assign tmp2122 = {const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0, const2121_0};
    assign tmp1502 = {temp_18[104], temp_18[105], temp_18[106], temp_18[107], temp_18[108], temp_18[109], temp_18[110], temp_18[111]};
    assign input_wire_9 = temp_31;
    assign tmp1998 = {tmp1997, tmp1805};
    assign tmp2419 = {const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0, const2418_0};
    assign tmp2657 = {temp_33[104], temp_33[105], temp_33[106], temp_33[107], temp_33[108], temp_33[109], temp_33[110], temp_33[111]};
    assign tmp2758 = tmp2754 ^ tmp2757;
    assign tmp388 = {const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0, const387_0};
    assign tmp1199 = {temp_13[48], temp_13[49], temp_13[50], temp_13[51], temp_13[52], temp_13[53], temp_13[54], temp_13[55]};
    assign tmp514 = tmp510 ^ tmp513;
        assign tmp1837 = mem_3[tmp1794];
        assign tmp995 = mem_4[tmp919];
    assign tmp1693 = {tmp1692, tmp1515};
    assign tmp1511 = {temp_18[32], temp_18[33], temp_18[34], temp_18[35], temp_18[36], temp_18[37], temp_18[38], temp_18[39]};
    assign tmp2581 = tmp2579 ^ tmp2580;
    assign temp_36 = new_10;
    assign tmp2213 = {tmp2212[0], tmp2212[1], tmp2212[2], tmp2212[3], tmp2212[4], tmp2212[5], tmp2212[6], tmp2212[7]};
    assign tmp640 = tmp700;
    assign tmp2793 = {tmp2792, tmp2677};
    assign tmp1718 = tmp1714 ^ tmp1717;
    assign tmp1195 = {temp_13[80], temp_13[81], temp_13[82], temp_13[83], temp_13[84], temp_13[85], temp_13[86], temp_13[87]};
    assign tmp2732 = {const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0, const2731_0};
    assign xor_w19 = tmp129;
    assign tmp2009 = {const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0, const2008_0};
        assign tmp1689 = mem_4[tmp1514];
    assign tmp1694 = tmp1690 ^ tmp1693;
        assign tmp396 = mem_3[tmp331];
    assign tmp1750 = tmp1766;
    assign tmp2681 = {temp_34[48], temp_34[49], temp_34[50], temp_34[51], temp_34[52], temp_34[53], temp_34[54], temp_34[55]};
        assign tmp1700 = mem_3[tmp1514];
        assign tmp1617 = mem_4[tmp1504];
        assign tmp2648 = mem_1[tmp2616];
    assign tmp428 = {const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0, const427_0};
    assign tmp366 = tmp362 ^ tmp365;
    assign tmp1526 = tmp1663;
    assign tmp1108 = tmp1104 ^ tmp1107;
    assign b3_w31 = tmp191;
        assign tmp2728 = mem_3[tmp2674];
    assign tmp1541 = {tmp1540, tmp1503};
    assign shifted_w3 = tmp13;
    assign tmp2816 = {const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0, const2815_0};
    assign tmp1913 = {const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0, const1912_0};
    assign new_9 = tmp2605;
    assign tmp416 = {const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0, const415_0};
    assign tmp2306 = {const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0, const2305_0};
    assign tmp2295 = {tmp2294, tmp2099};
    assign tmp2237 = {tmp2236[0], tmp2236[1], tmp2236[2], tmp2236[3], tmp2236[4], tmp2236[5], tmp2236[6], tmp2236[7]};
    assign tmp1530 = tmp1711;
    assign tmp2422 = {tmp2421[0], tmp2421[1], tmp2421[2], tmp2421[3], tmp2421[4], tmp2421[5], tmp2421[6], tmp2421[7]};
        assign tmp1934 = mem_4[tmp1803];
    assign tmp2796 = {const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0, const2795_0};
    assign tmp260 = {expanded_key[1280], expanded_key[1281], expanded_key[1282], expanded_key[1283], expanded_key[1284], expanded_key[1285], expanded_key[1286], expanded_key[1287], expanded_key[1288], expanded_key[1289], expanded_key[1290], expanded_key[1291], expanded_key[1292], expanded_key[1293], expanded_key[1294], expanded_key[1295], expanded_key[1296], expanded_key[1297], expanded_key[1298], expanded_key[1299], expanded_key[1300], expanded_key[1301], expanded_key[1302], expanded_key[1303], expanded_key[1304], expanded_key[1305], expanded_key[1306], expanded_key[1307], expanded_key[1308], expanded_key[1309], expanded_key[1310], expanded_key[1311], expanded_key[1312], expanded_key[1313], expanded_key[1314], expanded_key[1315], expanded_key[1316], expanded_key[1317], expanded_key[1318], expanded_key[1319], expanded_key[1320], expanded_key[1321], expanded_key[1322], expanded_key[1323], expanded_key[1324], expanded_key[1325], expanded_key[1326], expanded_key[1327], expanded_key[1328], expanded_key[1329], expanded_key[1330], expanded_key[1331], expanded_key[1332], expanded_key[1333], expanded_key[1334], expanded_key[1335], expanded_key[1336], expanded_key[1337], expanded_key[1338], expanded_key[1339], expanded_key[1340], expanded_key[1341], expanded_key[1342], expanded_key[1343], expanded_key[1344], expanded_key[1345], expanded_key[1346], expanded_key[1347], expanded_key[1348], expanded_key[1349], expanded_key[1350], expanded_key[1351], expanded_key[1352], expanded_key[1353], expanded_key[1354], expanded_key[1355], expanded_key[1356], expanded_key[1357], expanded_key[1358], expanded_key[1359], expanded_key[1360], expanded_key[1361], expanded_key[1362], expanded_key[1363], expanded_key[1364], expanded_key[1365], expanded_key[1366], expanded_key[1367], expanded_key[1368], expanded_key[1369], expanded_key[1370], expanded_key[1371], expanded_key[1372], expanded_key[1373], expanded_key[1374], expanded_key[1375], expanded_key[1376], expanded_key[1377], expanded_key[1378], expanded_key[1379], expanded_key[1380], expanded_key[1381], expanded_key[1382], expanded_key[1383], expanded_key[1384], expanded_key[1385], expanded_key[1386], expanded_key[1387], expanded_key[1388], expanded_key[1389], expanded_key[1390], expanded_key[1391], expanded_key[1392], expanded_key[1393], expanded_key[1394], expanded_key[1395], expanded_key[1396], expanded_key[1397], expanded_key[1398], expanded_key[1399], expanded_key[1400], expanded_key[1401], expanded_key[1402], expanded_key[1403], expanded_key[1404], expanded_key[1405], expanded_key[1406], expanded_key[1407]};
    assign tmp842 = {tmp841, tmp635};
    assign tmp932 = tmp981;
    assign tmp1406 = {tmp1405[0], tmp1405[1], tmp1405[2], tmp1405[3], tmp1405[4], tmp1405[5], tmp1405[6], tmp1405[7]};
    assign tmp434 = tmp432 ^ tmp433;
    assign tmp856 = {temp_8[56], temp_8[57], temp_8[58], temp_8[59], temp_8[60], temp_8[61], temp_8[62], temp_8[63]};
    assign tmp2337 = tmp2353;
    assign input_wire_8 = temp_27;
    assign tmp1566 = tmp1562 ^ tmp1565;
    assign tmp1672 = {const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0, const1671_0};
    assign tmp1283 = {const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0, const1282_0};
    assign tmp438 = tmp434 ^ tmp437;
        assign tmp2507 = mem_3[tmp2387];
    assign temp_19 = tmp1724;
        assign tmp68 = mem_1[b1_w11];
    assign tmp1756 = tmp1772;
    assign a2_w27 = tmp160;
    assign tmp1269 = tmp1265 ^ tmp1268;
        assign tmp224 = mem_2[const223_9];
    assign tmp1737 = {temp_20[40], temp_20[41], temp_20[42], temp_20[43], temp_20[44], temp_20[45], temp_20[46], temp_20[47]};
        assign tmp1300 = mem_4[tmp1213];
    assign tmp1438 = {temp_16[88], temp_16[89], temp_16[90], temp_16[91], temp_16[92], temp_16[93], temp_16[94], temp_16[95]};
    assign tmp2029 = {temp_24[48], temp_24[49], temp_24[50], temp_24[51], temp_24[52], temp_24[53], temp_24[54], temp_24[55]};
    assign b4_w3 = tmp17;
    assign tmp859 = {temp_8[32], temp_8[33], temp_8[34], temp_8[35], temp_8[36], temp_8[37], temp_8[38], temp_8[39]};
    assign tmp968 = tmp964 ^ tmp967;
    assign tmp1637 = {tmp1636, tmp1511};
    assign tmp2311 = {expanded_key[384], expanded_key[385], expanded_key[386], expanded_key[387], expanded_key[388], expanded_key[389], expanded_key[390], expanded_key[391], expanded_key[392], expanded_key[393], expanded_key[394], expanded_key[395], expanded_key[396], expanded_key[397], expanded_key[398], expanded_key[399], expanded_key[400], expanded_key[401], expanded_key[402], expanded_key[403], expanded_key[404], expanded_key[405], expanded_key[406], expanded_key[407], expanded_key[408], expanded_key[409], expanded_key[410], expanded_key[411], expanded_key[412], expanded_key[413], expanded_key[414], expanded_key[415], expanded_key[416], expanded_key[417], expanded_key[418], expanded_key[419], expanded_key[420], expanded_key[421], expanded_key[422], expanded_key[423], expanded_key[424], expanded_key[425], expanded_key[426], expanded_key[427], expanded_key[428], expanded_key[429], expanded_key[430], expanded_key[431], expanded_key[432], expanded_key[433], expanded_key[434], expanded_key[435], expanded_key[436], expanded_key[437], expanded_key[438], expanded_key[439], expanded_key[440], expanded_key[441], expanded_key[442], expanded_key[443], expanded_key[444], expanded_key[445], expanded_key[446], expanded_key[447], expanded_key[448], expanded_key[449], expanded_key[450], expanded_key[451], expanded_key[452], expanded_key[453], expanded_key[454], expanded_key[455], expanded_key[456], expanded_key[457], expanded_key[458], expanded_key[459], expanded_key[460], expanded_key[461], expanded_key[462], expanded_key[463], expanded_key[464], expanded_key[465], expanded_key[466], expanded_key[467], expanded_key[468], expanded_key[469], expanded_key[470], expanded_key[471], expanded_key[472], expanded_key[473], expanded_key[474], expanded_key[475], expanded_key[476], expanded_key[477], expanded_key[478], expanded_key[479], expanded_key[480], expanded_key[481], expanded_key[482], expanded_key[483], expanded_key[484], expanded_key[485], expanded_key[486], expanded_key[487], expanded_key[488], expanded_key[489], expanded_key[490], expanded_key[491], expanded_key[492], expanded_key[493], expanded_key[494], expanded_key[495], expanded_key[496], expanded_key[497], expanded_key[498], expanded_key[499], expanded_key[500], expanded_key[501], expanded_key[502], expanded_key[503], expanded_key[504], expanded_key[505], expanded_key[506], expanded_key[507], expanded_key[508], expanded_key[509], expanded_key[510], expanded_key[511]};
        assign tmp1557 = mem_4[tmp1503];
        assign tmp810 = mem_4[tmp635];
    assign tmp515 = {tmp514[0], tmp514[1], tmp514[2], tmp514[3], tmp514[4], tmp514[5], tmp514[6], tmp514[7]};
    assign c2_w31 = tmp194;
        assign tmp144 = mem_1[b2_w23];
    assign tmp1132 = tmp1128 ^ tmp1131;
    assign tmp204 = concat_w31 ^ substituted_w31;
    assign tmp1893 = {const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0, const1892_0};
    assign tmp722 = {tmp721, tmp625};
    assign tmp818 = {tmp817, tmp633};
    assign tmp282 = tmp298;
    assign tmp106 = tmp105 ^ tmp81;
    assign tmp724 = {tmp723[0], tmp723[1], tmp723[2], tmp723[3], tmp723[4], tmp723[5], tmp723[6], tmp723[7]};
    assign rc3_w35 = const226_0;
    assign tmp2673 = {temp_34[112], temp_34[113], temp_34[114], temp_34[115], temp_34[116], temp_34[117], temp_34[118], temp_34[119]};
    assign tmp506 = tmp504 ^ tmp505;
    assign tmp2159 = {tmp2158, tmp2087};
    assign tmp1094 = {const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0, const1093_0};
    assign tmp2160 = tmp2156 ^ tmp2159;
    assign rc4_w7 = const52_0;
        assign tmp958 = mem_3[tmp915];
    assign tmp567 = {temp_4[24], temp_4[25], temp_4[26], temp_4[27], temp_4[28], temp_4[29], temp_4[30], temp_4[31]};
    assign tmp1895 = tmp1891 ^ tmp1894;
    assign tmp1977 = {const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0, const1976_0};
    assign tmp1562 = tmp1558 ^ tmp1561;
        assign tmp602 = mem_1[tmp570];
    assign tmp2028 = {temp_24[56], temp_24[57], temp_24[58], temp_24[59], temp_24[60], temp_24[61], temp_24[62], temp_24[63]};
    assign tmp1525 = tmp1651;
    assign tmp1971 = tmp1969 ^ tmp1970;
    assign tmp2857 = {tmp2856, tmp2687};
    assign tmp976 = tmp972 ^ tmp975;
    assign tmp662 = {tmp661, tmp624};
    assign tmp2129 = {tmp2128[0], tmp2128[1], tmp2128[2], tmp2128[3], tmp2128[4], tmp2128[5], tmp2128[6], tmp2128[7]};
    assign tmp2254 = {const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0, const2253_0};
    assign tmp2622 = tmp2638;
    assign tmp264 = {new_state[104], new_state[105], new_state[106], new_state[107], new_state[108], new_state[109], new_state[110], new_state[111]};
    assign tmp1249 = tmp1245 ^ tmp1248;
    assign tmp208 = tmp207 ^ tmp183;
    assign tmp1150 = {temp_12[48], temp_12[49], temp_12[50], temp_12[51], temp_12[52], temp_12[53], temp_12[54], temp_12[55]};
    assign b1_w23 = tmp139;
    assign tmp2413 = tmp2411 ^ tmp2412;
        assign tmp170 = mem_1[b3_w27];
    assign tmp466 = tmp462 ^ tmp465;
    assign tmp733 = {const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0, const732_0};
    assign tmp651 = tmp832;
        assign tmp1182 = mem_1[tmp1150];
    assign tmp479 = {tmp478[0], tmp478[1], tmp478[2], tmp478[3], tmp478[4], tmp478[5], tmp478[6], tmp478[7]};
        assign tmp1054 = mem_3[tmp923];
    assign tmp1567 = {tmp1566[0], tmp1566[1], tmp1566[2], tmp1566[3], tmp1566[4], tmp1566[5], tmp1566[6], tmp1566[7]};
    assign tmp22 = {c1_w3, c2_w3, c3_w3, c4_w3};
    assign tmp2318 = {temp_28[80], temp_28[81], temp_28[82], temp_28[83], temp_28[84], temp_28[85], temp_28[86], temp_28[87]};
    assign tmp1589 = {tmp1588, tmp1507};
        assign tmp587 = mem_1[tmp555];
        assign tmp798 = mem_4[tmp634];
    assign tmp478 = tmp474 ^ tmp477;
        assign tmp1544 = mem_3[tmp1501];
    assign tmp2073 = {temp_25[88], temp_25[89], temp_25[90], temp_25[91], temp_25[92], temp_25[93], temp_25[94], temp_25[95]};
    assign tmp2493 = tmp2489 ^ tmp2492;
        assign tmp1909 = mem_3[tmp1800];
    assign tmp1449 = {temp_16[0], temp_16[1], temp_16[2], temp_16[3], temp_16[4], temp_16[5], temp_16[6], temp_16[7]};
        assign tmp2119 = mem_4[tmp2087];
    assign tmp140 = {shifted_w23[16], shifted_w23[17], shifted_w23[18], shifted_w23[19], shifted_w23[20], shifted_w23[21], shifted_w23[22], shifted_w23[23]};
    assign rc2_w27 = const175_0;
    assign tmp1161 = tmp1177;
    assign tmp2290 = {const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0, const2289_0};
    assign tmp550 = tmp546 ^ tmp549;
    assign tmp2343 = tmp2359;
    assign tmp646 = tmp772;
    assign tmp2709 = {tmp2708, tmp2674};
    assign temp_37 = tmp2947;
        assign tmp749 = mem_3[tmp629];
    assign tmp240 = {shifted_w39[16], shifted_w39[17], shifted_w39[18], shifted_w39[19], shifted_w39[20], shifted_w39[21], shifted_w39[22], shifted_w39[23]};
    assign tmp1704 = {const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0, const1703_0};
    assign tmp131 = tmp130 ^ tmp106;
    assign tmp2404 = tmp2530;
    assign tmp2476 = {tmp2475, tmp2386};
    assign tmp645 = tmp760;
    assign tmp1465 = tmp1481;
    assign tmp2757 = {tmp2756, tmp2678};
    assign tmp617 = {temp_5[16], temp_5[17], temp_5[18], temp_5[19], temp_5[20], temp_5[21], temp_5[22], temp_5[23]};
    assign tmp1309 = tmp1305 ^ tmp1308;
    assign tmp903 = {temp_9[72], temp_9[73], temp_9[74], temp_9[75], temp_9[76], temp_9[77], temp_9[78], temp_9[79]};
    assign w7 = tmp33;
    assign tmp2420 = {tmp2419, tmp2382};
    assign b3_w7 = tmp41;
        assign tmp2353 = mem_1[tmp2321];
    assign tmp289 = tmp305;
    assign temp_27 = tmp2310;
        assign tmp397 = mem_4[tmp328];
    assign tmp852 = {temp_8[88], temp_8[89], temp_8[90], temp_8[91], temp_8[92], temp_8[93], temp_8[94], temp_8[95]};
    assign input_wire_6 = temp_19;
    assign tmp2736 = {const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0, const2735_0};
    assign tmp2140 = tmp2136 ^ tmp2139;
    assign tmp1382 = {tmp1381[0], tmp1381[1], tmp1381[2], tmp1381[3], tmp1381[4], tmp1381[5], tmp1381[6], tmp1381[7]};
    assign new_11 = tmp2966;
    assign tmp1792 = {tmp1776, tmp1781, tmp1786, tmp1791, tmp1780, tmp1785, tmp1790, tmp1779, tmp1784, tmp1789, tmp1778, tmp1783, tmp1788, tmp1777, tmp1782, tmp1787};
    assign tmp2677 = {temp_34[80], temp_34[81], temp_34[82], temp_34[83], temp_34[84], temp_34[85], temp_34[86], temp_34[87]};
    assign tmp2790 = tmp2788 ^ tmp2789;
    assign tmp2666 = {temp_33[32], temp_33[33], temp_33[34], temp_33[35], temp_33[36], temp_33[37], temp_33[38], temp_33[39]};
    assign tmp2437 = tmp2435 ^ tmp2436;
    assign tmp2176 = tmp2172 ^ tmp2175;
        assign tmp666 = mem_4[tmp623];
    assign tmp1951 = tmp1947 ^ tmp1950;
    assign tmp2452 = {tmp2451, tmp2380};
    assign tmp1795 = {temp_22[104], temp_22[105], temp_22[106], temp_22[107], temp_22[108], temp_22[109], temp_22[110], temp_22[111]};
    assign tmp1068 = tmp1066 ^ tmp1067;
    assign tmp192 = {shifted_w31[0], shifted_w31[1], shifted_w31[2], shifted_w31[3], shifted_w31[4], shifted_w31[5], shifted_w31[6], shifted_w31[7]};
    assign tmp2847 = {tmp2846[0], tmp2846[1], tmp2846[2], tmp2846[3], tmp2846[4], tmp2846[5], tmp2846[6], tmp2846[7]};
    assign tmp1819 = tmp1956;
    assign tmp613 = {temp_5[48], temp_5[49], temp_5[50], temp_5[51], temp_5[52], temp_5[53], temp_5[54], temp_5[55]};
    assign tmp1486 = {temp_17[96], temp_17[97], temp_17[98], temp_17[99], temp_17[100], temp_17[101], temp_17[102], temp_17[103]};
    assign tmp783 = tmp779 ^ tmp782;
    assign tmp1087 = {tmp1086, tmp924};
    assign tmp1307 = {const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0, const1306_0};
    assign tmp1776 = {temp_21[120], temp_21[121], temp_21[122], temp_21[123], temp_21[124], temp_21[125], temp_21[126], temp_21[127]};
    assign tmp133 = tmp132 ^ tmp108;
    assign tmp2283 = {tmp2282, tmp2098};
    assign tmp239 = {shifted_w39[24], shifted_w39[25], shifted_w39[26], shifted_w39[27], shifted_w39[28], shifted_w39[29], shifted_w39[30], shifted_w39[31]};
    assign tmp866 = tmp882;
    assign tmp2805 = {tmp2804, tmp2682};
    assign b2_w27 = tmp165;
    assign tmp2835 = {tmp2834[0], tmp2834[1], tmp2834[2], tmp2834[3], tmp2834[4], tmp2834[5], tmp2834[6], tmp2834[7]};
    assign tmp980 = tmp976 ^ tmp979;
    assign tmp1445 = {temp_16[32], temp_16[33], temp_16[34], temp_16[35], temp_16[36], temp_16[37], temp_16[38], temp_16[39]};
    assign tmp860 = {temp_8[24], temp_8[25], temp_8[26], temp_8[27], temp_8[28], temp_8[29], temp_8[30], temp_8[31]};
        assign tmp597 = mem_1[tmp565];
    assign tmp2036 = tmp2052;
    assign tmp2247 = {tmp2246, tmp2095};
        assign tmp2944 = mem_1[tmp2912];
    assign b1_w15 = tmp89;
    assign tmp1757 = tmp1773;
    assign tmp1917 = {const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0, const1916_0};
    assign tmp2882 = tmp2878 ^ tmp2881;
    assign tmp182 = tmp181 ^ tmp157;
    assign tmp2096 = {temp_26[40], temp_26[41], temp_26[42], temp_26[43], temp_26[44], temp_26[45], temp_26[46], temp_26[47]};
    assign tmp2128 = tmp2124 ^ tmp2127;
        assign tmp243 = mem_1[b1_w39];
    assign tmp937 = tmp1041;
    assign tmp2021 = {temp_24[112], temp_24[113], temp_24[114], temp_24[115], temp_24[116], temp_24[117], temp_24[118], temp_24[119]};
        assign tmp69 = mem_1[b2_w11];
    assign tmp1310 = {tmp1309[0], tmp1309[1], tmp1309[2], tmp1309[3], tmp1309[4], tmp1309[5], tmp1309[6], tmp1309[7]};
        assign tmp821 = mem_3[tmp635];
    assign tmp1706 = tmp1702 ^ tmp1705;
    assign tmp1510 = {temp_18[40], temp_18[41], temp_18[42], temp_18[43], temp_18[44], temp_18[45], temp_18[46], temp_18[47]};
        assign tmp2472 = mem_4[tmp2385];
        assign tmp971 = mem_4[tmp917];
    assign tmp2477 = tmp2473 ^ tmp2476;
        assign tmp297 = mem_1[tmp265];
        assign tmp1372 = mem_4[tmp1215];
    assign tmp2635 = tmp2651;
        assign tmp420 = mem_3[tmp333];
    assign tmp2204 = tmp2202 ^ tmp2203;
    assign tmp931 = tmp969;
    assign tmp936 = tmp1029;
    assign tmp512 = {const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0, const511_0};
    assign tmp115 = {shifted_w19[16], shifted_w19[17], shifted_w19[18], shifted_w19[19], shifted_w19[20], shifted_w19[21], shifted_w19[22], shifted_w19[23]};
    assign tmp1169 = tmp1185;
    assign rc3_w31 = const201_0;
    assign tmp657 = {const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0, const656_0};
    assign tmp1927 = tmp1923 ^ tmp1926;
        assign tmp946 = mem_3[tmp914];
        assign tmp1862 = mem_4[tmp1793];
    assign tmp1938 = {tmp1937, tmp1804};
    assign b2_w3 = tmp15;
    assign tmp2606 = {temp_32[120], temp_32[121], temp_32[122], temp_32[123], temp_32[124], temp_32[125], temp_32[126], temp_32[127]};
    assign tmp2954 = {temp_37[72], temp_37[73], temp_37[74], temp_37[75], temp_37[76], temp_37[77], temp_37[78], temp_37[79]};
        assign tmp762 = mem_4[tmp631];
    assign a4_w27 = tmp162;
    assign tmp1096 = tmp1092 ^ tmp1095;
        assign tmp1957 = mem_3[tmp1804];
    assign tmp1434 = {temp_16[120], temp_16[121], temp_16[122], temp_16[123], temp_16[124], temp_16[125], temp_16[126], temp_16[127]};
    assign rc1_w35 = tmp224;
    assign tmp614 = {temp_5[40], temp_5[41], temp_5[42], temp_5[43], temp_5[44], temp_5[45], temp_5[46], temp_5[47]};
    assign tmp1999 = tmp1995 ^ tmp1998;
    assign tmp448 = {const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0, const447_0};
    assign tmp1965 = {const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0, const1964_0};
    assign tmp326 = {temp_1[0], temp_1[1], temp_1[2], temp_1[3], temp_1[4], temp_1[5], temp_1[6], temp_1[7]};
        assign tmp1768 = mem_1[tmp1736];
    assign input_wire_5 = temp_15;
    assign tmp2230 = {const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0, const2229_0};
    assign b1_w3 = tmp14;
    assign tmp553 = {expanded_key[1152], expanded_key[1153], expanded_key[1154], expanded_key[1155], expanded_key[1156], expanded_key[1157], expanded_key[1158], expanded_key[1159], expanded_key[1160], expanded_key[1161], expanded_key[1162], expanded_key[1163], expanded_key[1164], expanded_key[1165], expanded_key[1166], expanded_key[1167], expanded_key[1168], expanded_key[1169], expanded_key[1170], expanded_key[1171], expanded_key[1172], expanded_key[1173], expanded_key[1174], expanded_key[1175], expanded_key[1176], expanded_key[1177], expanded_key[1178], expanded_key[1179], expanded_key[1180], expanded_key[1181], expanded_key[1182], expanded_key[1183], expanded_key[1184], expanded_key[1185], expanded_key[1186], expanded_key[1187], expanded_key[1188], expanded_key[1189], expanded_key[1190], expanded_key[1191], expanded_key[1192], expanded_key[1193], expanded_key[1194], expanded_key[1195], expanded_key[1196], expanded_key[1197], expanded_key[1198], expanded_key[1199], expanded_key[1200], expanded_key[1201], expanded_key[1202], expanded_key[1203], expanded_key[1204], expanded_key[1205], expanded_key[1206], expanded_key[1207], expanded_key[1208], expanded_key[1209], expanded_key[1210], expanded_key[1211], expanded_key[1212], expanded_key[1213], expanded_key[1214], expanded_key[1215], expanded_key[1216], expanded_key[1217], expanded_key[1218], expanded_key[1219], expanded_key[1220], expanded_key[1221], expanded_key[1222], expanded_key[1223], expanded_key[1224], expanded_key[1225], expanded_key[1226], expanded_key[1227], expanded_key[1228], expanded_key[1229], expanded_key[1230], expanded_key[1231], expanded_key[1232], expanded_key[1233], expanded_key[1234], expanded_key[1235], expanded_key[1236], expanded_key[1237], expanded_key[1238], expanded_key[1239], expanded_key[1240], expanded_key[1241], expanded_key[1242], expanded_key[1243], expanded_key[1244], expanded_key[1245], expanded_key[1246], expanded_key[1247], expanded_key[1248], expanded_key[1249], expanded_key[1250], expanded_key[1251], expanded_key[1252], expanded_key[1253], expanded_key[1254], expanded_key[1255], expanded_key[1256], expanded_key[1257], expanded_key[1258], expanded_key[1259], expanded_key[1260], expanded_key[1261], expanded_key[1262], expanded_key[1263], expanded_key[1264], expanded_key[1265], expanded_key[1266], expanded_key[1267], expanded_key[1268], expanded_key[1269], expanded_key[1270], expanded_key[1271], expanded_key[1272], expanded_key[1273], expanded_key[1274], expanded_key[1275], expanded_key[1276], expanded_key[1277], expanded_key[1278], expanded_key[1279]};
    assign tmp2470 = {tmp2469[0], tmp2469[1], tmp2469[2], tmp2469[3], tmp2469[4], tmp2469[5], tmp2469[6], tmp2469[7]};
    assign tmp1431 = {tmp1223, tmp1224, tmp1225, tmp1226, tmp1227, tmp1228, tmp1229, tmp1230, tmp1231, tmp1232, tmp1233, tmp1234, tmp1235, tmp1236, tmp1237, tmp1238};
    assign tmp2631 = tmp2647;
        assign tmp1605 = mem_4[tmp1507];
    assign tmp325 = {temp_1[8], temp_1[9], temp_1[10], temp_1[11], temp_1[12], temp_1[13], temp_1[14], temp_1[15]};
    assign b1_w11 = tmp64;
    assign tmp545 = {tmp544, tmp341};
    assign tmp2660 = {temp_33[80], temp_33[81], temp_33[82], temp_33[83], temp_33[84], temp_33[85], temp_33[86], temp_33[87]};
    assign concat_w3 = tmp28;
    assign tmp15 = {shifted_w3[16], shifted_w3[17], shifted_w3[18], shifted_w3[19], shifted_w3[20], shifted_w3[21], shifted_w3[22], shifted_w3[23]};
    assign tmp580 = tmp596;
    assign tmp1058 = {const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0, const1057_0};
    assign tmp2821 = {tmp2820, tmp2680};
    assign tmp1645 = {tmp1644, tmp1511};
    assign a2_w35 = tmp210;
    assign tmp1843 = tmp1839 ^ tmp1842;
    assign input_wire_1 = aes_plaintext;
    assign tmp429 = {tmp428, tmp332};
    assign tmp572 = tmp588;
    assign tmp925 = {temp_10[32], temp_10[33], temp_10[34], temp_10[35], temp_10[36], temp_10[37], temp_10[38], temp_10[39]};
        assign tmp385 = mem_4[tmp331];
    assign tmp1986 = {tmp1985, tmp1808};
        assign tmp219 = mem_1[b2_w35];
    assign c3_w3 = tmp20;
    assign tmp634 = {temp_6[16], temp_6[17], temp_6[18], temp_6[19], temp_6[20], temp_6[21], temp_6[22], temp_6[23]};
    assign tmp154 = concat_w23 ^ substituted_w23;
    assign tmp2599 = {const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0, const2598_0};
    assign tmp709 = {const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0, const708_0};
    assign tmp1882 = {tmp1881, tmp1800};
    assign tmp1968 = {tmp1967[0], tmp1967[1], tmp1967[2], tmp1967[3], tmp1967[4], tmp1967[5], tmp1967[6], tmp1967[7]};
    assign tmp2683 = {temp_34[32], temp_34[33], temp_34[34], temp_34[35], temp_34[36], temp_34[37], temp_34[38], temp_34[39]};
    assign tmp1011 = {tmp1010, tmp921};
    assign tmp1106 = {const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0, const1105_0};
    assign tmp2702 = tmp2883;
    assign tmp2818 = tmp2814 ^ tmp2817;
    assign tmp36 = {w7[8], w7[9], w7[10], w7[11], w7[12], w7[13], w7[14], w7[15]};
    assign temp_2 = tmp327;
    assign tmp485 = {tmp484, tmp336};
    assign tmp942 = tmp1101;
    assign tmp72 = {c1_w11, c2_w11, c3_w11, c4_w11};
    assign tmp39 = {shifted_w7[24], shifted_w7[25], shifted_w7[26], shifted_w7[27], shifted_w7[28], shifted_w7[29], shifted_w7[30], shifted_w7[31]};
        assign tmp469 = mem_4[tmp338];
    assign tmp817 = {const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0, const816_0};
    assign tmp1214 = {temp_14[64], temp_14[65], temp_14[66], temp_14[67], temp_14[68], temp_14[69], temp_14[70], temp_14[71]};
    assign tmp2920 = tmp2936;
    assign tmp2076 = {temp_25[64], temp_25[65], temp_25[66], temp_25[67], temp_25[68], temp_25[69], temp_25[70], temp_25[71]};
        assign tmp2943 = mem_1[tmp2911];
    assign tmp1225 = tmp1274;
    assign tmp778 = {tmp777, tmp629};
    assign tmp1156 = {temp_12[0], temp_12[1], temp_12[2], temp_12[3], temp_12[4], temp_12[5], temp_12[6], temp_12[7]};
        assign tmp1873 = mem_3[tmp1797];
    assign xor_w11 = tmp79;
    assign xor_w27 = tmp179;
    assign tmp1076 = tmp1072 ^ tmp1075;
        assign tmp2352 = mem_1[tmp2320];
    assign tmp2619 = {temp_32[16], temp_32[17], temp_32[18], temp_32[19], temp_32[20], temp_32[21], temp_32[22], temp_32[23]};
    assign tmp2722 = tmp2718 ^ tmp2721;
    assign tmp1256 = {tmp1255, tmp1210};
    assign tmp851 = {temp_8[96], temp_8[97], temp_8[98], temp_8[99], temp_8[100], temp_8[101], temp_8[102], temp_8[103]};
        assign tmp2298 = mem_3[tmp2101];
        assign tmp2052 = mem_1[tmp2020];
        assign tmp725 = mem_3[tmp627];
        assign tmp2646 = mem_1[tmp2614];
        assign tmp2651 = mem_1[tmp2619];
    assign tmp2698 = tmp2835;
    assign tmp1709 = {tmp1708, tmp1513};
        assign tmp2360 = mem_1[tmp2328];
    assign tmp1453 = tmp1469;
    assign tmp2210 = {const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0, const2209_0};
    assign tmp1633 = {tmp1632, tmp1510};
    assign tmp2141 = {tmp2140[0], tmp2140[1], tmp2140[2], tmp2140[3], tmp2140[4], tmp2140[5], tmp2140[6], tmp2140[7]};
        assign tmp598 = mem_1[tmp566];
    assign tmp1429 = tmp1425 ^ tmp1428;
        assign tmp887 = mem_1[tmp855];
    assign tmp2002 = {tmp2001, tmp1806};
    assign tmp1531 = tmp1723;
    assign tmp2249 = {tmp2248[0], tmp2248[1], tmp2248[2], tmp2248[3], tmp2248[4], tmp2248[5], tmp2248[6], tmp2248[7]};
    assign tmp1889 = {const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0, const1888_0};
    assign tmp899 = {temp_9[104], temp_9[105], temp_9[106], temp_9[107], temp_9[108], temp_9[109], temp_9[110], temp_9[111]};
    assign tmp1341 = tmp1337 ^ tmp1340;
    assign tmp2082 = {temp_25[16], temp_25[17], temp_25[18], temp_25[19], temp_25[20], temp_25[21], temp_25[22], temp_25[23]};
    assign tmp2901 = {temp_36[104], temp_36[105], temp_36[106], temp_36[107], temp_36[108], temp_36[109], temp_36[110], temp_36[111]};
    assign tmp530 = tmp528 ^ tmp529;
    assign tmp1914 = {tmp1913, tmp1798};
        assign tmp2239 = mem_4[tmp2097];
    assign tmp1809 = tmp1836;
    assign tmp2734 = tmp2730 ^ tmp2733;
    assign tmp1735 = {temp_20[56], temp_20[57], temp_20[58], temp_20[59], temp_20[60], temp_20[61], temp_20[62], temp_20[63]};
    assign tmp1203 = {temp_13[16], temp_13[17], temp_13[18], temp_13[19], temp_13[20], temp_13[21], temp_13[22], temp_13[23]};
        assign tmp517 = mem_4[tmp342];
    assign tmp2817 = {tmp2816, tmp2683};
    assign tmp2396 = tmp2434;
        assign tmp2191 = mem_4[tmp2093];
    assign tmp1781 = {temp_21[80], temp_21[81], temp_21[82], temp_21[83], temp_21[84], temp_21[85], temp_21[86], temp_21[87]};
    assign tmp939 = tmp1065;
        assign tmp2940 = mem_1[tmp2908];
    assign tmp2671 = {tmp2655, tmp2660, tmp2665, tmp2670, tmp2659, tmp2664, tmp2669, tmp2658, tmp2663, tmp2668, tmp2657, tmp2662, tmp2667, tmp2656, tmp2661, tmp2666};
    assign a4_w23 = tmp137;
    assign tmp2409 = tmp2590;
    assign tmp736 = {tmp735[0], tmp735[1], tmp735[2], tmp735[3], tmp735[4], tmp735[5], tmp735[6], tmp735[7]};
    assign substituted_w23 = tmp147;
    assign tmp2910 = {temp_36[32], temp_36[33], temp_36[34], temp_36[35], temp_36[36], temp_36[37], temp_36[38], temp_36[39]};
    assign a2_w39 = tmp235;
    assign tmp1829 = {const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0, const1828_0};
    assign tmp424 = {const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0, const423_0};
    assign xor_w35 = tmp229;
    assign tmp338 = {temp_2[40], temp_2[41], temp_2[42], temp_2[43], temp_2[44], temp_2[45], temp_2[46], temp_2[47]};
    assign tmp2593 = tmp2591 ^ tmp2592;
    assign tmp1118 = {const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0, const1117_0};
    assign tmp455 = {tmp454[0], tmp454[1], tmp454[2], tmp454[3], tmp454[4], tmp454[5], tmp454[6], tmp454[7]};
    assign tmp1357 = tmp1353 ^ tmp1356;
    assign tmp1447 = {temp_16[16], temp_16[17], temp_16[18], temp_16[19], temp_16[20], temp_16[21], temp_16[22], temp_16[23]};
        assign tmp2591 = mem_3[tmp2394];
    assign tmp898 = {temp_9[112], temp_9[113], temp_9[114], temp_9[115], temp_9[116], temp_9[117], temp_9[118], temp_9[119]};
    assign tmp1923 = tmp1921 ^ tmp1922;
    assign tmp2451 = {const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0, const2450_0};
    assign tmp839 = tmp835 ^ tmp838;
    assign tmp1015 = {tmp1014, tmp918};
        assign tmp1179 = mem_1[tmp1147];
    assign tmp912 = {temp_9[0], temp_9[1], temp_9[2], temp_9[3], temp_9[4], temp_9[5], temp_9[6], temp_9[7]};
    assign tmp2225 = {tmp2224[0], tmp2224[1], tmp2224[2], tmp2224[3], tmp2224[4], tmp2224[5], tmp2224[6], tmp2224[7]};
        assign tmp2652 = mem_1[tmp2620];
    assign tmp354 = tmp491;
    assign tmp1418 = {tmp1417[0], tmp1417[1], tmp1417[2], tmp1417[3], tmp1417[4], tmp1417[5], tmp1417[6], tmp1417[7]};
    assign tmp1749 = tmp1765;
    assign tmp659 = tmp655 ^ tmp658;
    assign tmp2708 = {const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0, const2707_0};
        assign tmp726 = mem_4[tmp628];
    assign tmp987 = {tmp986, tmp915};
    assign tmp323 = {temp_1[24], temp_1[25], temp_1[26], temp_1[27], temp_1[28], temp_1[29], temp_1[30], temp_1[31]};
    assign tmp5 = {aes_key[96], aes_key[97], aes_key[98], aes_key[99], aes_key[100], aes_key[101], aes_key[102], aes_key[103], aes_key[104], aes_key[105], aes_key[106], aes_key[107], aes_key[108], aes_key[109], aes_key[110], aes_key[111], aes_key[112], aes_key[113], aes_key[114], aes_key[115], aes_key[116], aes_key[117], aes_key[118], aes_key[119], aes_key[120], aes_key[121], aes_key[122], aes_key[123], aes_key[124], aes_key[125], aes_key[126], aes_key[127]};
    assign tmp2223 = {tmp2222, tmp2097};
    assign tmp674 = {tmp673, tmp621};
    assign tmp2317 = {temp_28[88], temp_28[89], temp_28[90], temp_28[91], temp_28[92], temp_28[93], temp_28[94], temp_28[95]};
    assign tmp2284 = tmp2280 ^ tmp2283;
        assign tmp2227 = mem_4[tmp2096];
    assign tmp1806 = {temp_22[16], temp_22[17], temp_22[18], temp_22[19], temp_22[20], temp_22[21], temp_22[22], temp_22[23]};
    assign tmp2457 = tmp2453 ^ tmp2456;
    assign tmp2770 = tmp2766 ^ tmp2769;
        assign tmp2059 = mem_1[tmp2027];
        assign tmp1604 = mem_3[tmp1506];
    assign tmp336 = {temp_2[56], temp_2[57], temp_2[58], temp_2[59], temp_2[60], temp_2[61], temp_2[62], temp_2[63]};
        assign tmp1712 = mem_3[tmp1515];
    assign tmp1942 = {tmp1941, tmp1801};
    assign tmp875 = tmp891;
    assign tmp566 = {temp_4[32], temp_4[33], temp_4[34], temp_4[35], temp_4[36], temp_4[37], temp_4[38], temp_4[39]};
    assign tmp355 = tmp503;
    assign tmp1869 = {const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0, const1868_0};
        assign tmp2776 = mem_3[tmp2678];
    assign tmp1430 = {tmp1429[0], tmp1429[1], tmp1429[2], tmp1429[3], tmp1429[4], tmp1429[5], tmp1429[6], tmp1429[7]};
    assign tmp698 = {tmp697, tmp623};
    assign tmp2439 = {const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0, const2438_0};
        assign tmp457 = mem_4[tmp337];
    assign tmp1705 = {tmp1704, tmp1512};
    assign tmp2334 = tmp2350;
    assign tmp1157 = tmp1173;
    assign tmp80 = tmp55 ^ xor_w11;
    assign tmp1454 = tmp1470;
    assign tmp383 = {tmp382[0], tmp382[1], tmp382[2], tmp382[3], tmp382[4], tmp382[5], tmp382[6], tmp382[7]};
    assign tmp1305 = tmp1301 ^ tmp1304;
    assign tmp37 = {w7[0], w7[1], w7[2], w7[3], w7[4], w7[5], w7[6], w7[7]};
    assign w2 = tmp7;
        assign tmp2650 = mem_1[tmp2618];
    assign tmp544 = {const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0, const543_0};
    assign tmp2890 = tmp2886 ^ tmp2889;
    assign tmp2785 = {tmp2784, tmp2677};
    assign tmp896 = {tmp864, tmp865, tmp866, tmp867, tmp868, tmp869, tmp870, tmp871, tmp872, tmp873, tmp874, tmp875, tmp876, tmp877, tmp878, tmp879};
    assign tmp872 = tmp888;
    assign tmp2316 = {temp_28[96], temp_28[97], temp_28[98], temp_28[99], temp_28[100], temp_28[101], temp_28[102], temp_28[103]};
        assign tmp595 = mem_1[tmp563];
        assign tmp1770 = mem_1[tmp1738];
        assign tmp2592 = mem_4[tmp2391];
    assign tmp2896 = {tmp2688, tmp2689, tmp2690, tmp2691, tmp2692, tmp2693, tmp2694, tmp2695, tmp2696, tmp2697, tmp2698, tmp2699, tmp2700, tmp2701, tmp2702, tmp2703};
        assign tmp2532 = mem_4[tmp2390];
        assign tmp2508 = mem_4[tmp2388];
    assign tmp167 = {shifted_w27[0], shifted_w27[1], shifted_w27[2], shifted_w27[3], shifted_w27[4], shifted_w27[5], shifted_w27[6], shifted_w27[7]};
    assign tmp2074 = {temp_25[80], temp_25[81], temp_25[82], temp_25[83], temp_25[84], temp_25[85], temp_25[86], temp_25[87]};
    assign tmp2077 = {temp_25[56], temp_25[57], temp_25[58], temp_25[59], temp_25[60], temp_25[61], temp_25[62], temp_25[63]};
    assign c3_w19 = tmp120;
    assign tmp2078 = {temp_25[48], temp_25[49], temp_25[50], temp_25[51], temp_25[52], temp_25[53], temp_25[54], temp_25[55]};
    assign a1_w35 = tmp209;
        assign tmp361 = mem_4[tmp329];
    assign tmp2750 = tmp2746 ^ tmp2749;
    assign tmp1721 = {tmp1720, tmp1514};
        assign tmp1240 = mem_4[tmp1208];
    assign b4_w15 = tmp92;
    assign tmp255 = tmp230 ^ xor_w39;
    assign tmp2492 = {tmp2491, tmp2384};
        assign tmp408 = mem_3[tmp332];
    assign tmp1333 = tmp1329 ^ tmp1332;
    assign w0 = tmp5;
    assign tmp1344 = {tmp1343, tmp1218};
    assign tmp2443 = {const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0, const2442_0};
    assign tmp2222 = {const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0, const2221_0};
    assign tmp2187 = {tmp2186, tmp2090};
    assign tmp2297 = {tmp2296[0], tmp2296[1], tmp2296[2], tmp2296[3], tmp2296[4], tmp2296[5], tmp2296[6], tmp2296[7]};
        assign tmp1970 = mem_4[tmp1806];
    assign tmp772 = {tmp771[0], tmp771[1], tmp771[2], tmp771[3], tmp771[4], tmp771[5], tmp771[6], tmp771[7]};
    assign tmp2256 = tmp2252 ^ tmp2255;
    assign tmp2956 = {temp_37[56], temp_37[57], temp_37[58], temp_37[59], temp_37[60], temp_37[61], temp_37[62], temp_37[63]};
    assign tmp2900 = {temp_36[112], temp_36[113], temp_36[114], temp_36[115], temp_36[116], temp_36[117], temp_36[118], temp_36[119]};
    assign temp_25 = tmp2068;
    assign tmp1448 = {temp_16[8], temp_16[9], temp_16[10], temp_16[11], temp_16[12], temp_16[13], temp_16[14], temp_16[15]};
    assign tmp410 = tmp408 ^ tmp409;
        assign tmp2849 = mem_4[tmp2685];
    assign tmp316 = {temp_1[80], temp_1[81], temp_1[82], temp_1[83], temp_1[84], temp_1[85], temp_1[86], temp_1[87]};
    assign tmp402 = tmp398 ^ tmp401;
    assign tmp2458 = {tmp2457[0], tmp2457[1], tmp2457[2], tmp2457[3], tmp2457[4], tmp2457[5], tmp2457[6], tmp2457[7]};
    assign a4_w31 = tmp187;
    assign tmp1024 = tmp1020 ^ tmp1023;
        assign tmp689 = mem_3[tmp624];
    assign tmp1008 = tmp1006 ^ tmp1007;
        assign tmp2931 = mem_1[tmp2899];
    assign tmp1620 = {const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0, const1619_0};
    assign tmp1193 = {temp_13[96], temp_13[97], temp_13[98], temp_13[99], temp_13[100], temp_13[101], temp_13[102], temp_13[103]};
    assign tmp1650 = tmp1646 ^ tmp1649;
    assign tmp928 = {temp_10[8], temp_10[9], temp_10[10], temp_10[11], temp_10[12], temp_10[13], temp_10[14], temp_10[15]};
    assign tmp2878 = tmp2874 ^ tmp2877;
        assign tmp1764 = mem_1[tmp1732];
    assign tmp1381 = tmp1377 ^ tmp1380;
    assign tmp1901 = {const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0, const1900_0};
    assign tmp559 = {temp_4[88], temp_4[89], temp_4[90], temp_4[91], temp_4[92], temp_4[93], temp_4[94], temp_4[95]};
    assign tmp2808 = {const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0, const2807_0};
    assign tmp789 = {const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0, const788_0};
    assign tmp948 = tmp946 ^ tmp947;
    assign tmp1902 = {tmp1901, tmp1797};
    assign tmp907 = {temp_9[40], temp_9[41], temp_9[42], temp_9[43], temp_9[44], temp_9[45], temp_9[46], temp_9[47]};
        assign tmp44 = mem_1[b2_w7];
    assign tmp1241 = tmp1239 ^ tmp1240;
    assign temp_1 = tmp310;
    assign tmp1500 = {temp_18[120], temp_18[121], temp_18[122], temp_18[123], temp_18[124], temp_18[125], temp_18[126], temp_18[127]};
    assign tmp1301 = tmp1299 ^ tmp1300;
    assign tmp2280 = tmp2276 ^ tmp2279;
    assign tmp1801 = {temp_22[56], temp_22[57], temp_22[58], temp_22[59], temp_22[60], temp_22[61], temp_22[62], temp_22[63]};
    assign tmp2892 = {const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0, const2891_0};
    assign tmp2503 = {const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0, const2502_0};
    assign temp_22 = tmp1792;
        assign tmp1115 = mem_4[tmp929];
    assign tmp718 = {tmp717, tmp628};
    assign tmp2889 = {tmp2888, tmp2685};
    assign tmp29 = concat_w3 ^ substituted_w3;
    assign substituted_w15 = tmp97;
    assign tmp1046 = {const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0, const1045_0};
        assign tmp2556 = mem_4[tmp2392];
    assign tmp2588 = {tmp2587, tmp2392};
    assign tmp2124 = tmp2120 ^ tmp2123;
    assign tmp835 = tmp833 ^ tmp834;
    assign tmp1002 = {const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0, const1001_0};
    assign tmp2907 = {temp_36[56], temp_36[57], temp_36[58], temp_36[59], temp_36[60], temp_36[61], temp_36[62], temp_36[63]};
    assign rc4_w19 = const127_0;
    assign tmp1834 = {tmp1833, tmp1796};
        assign tmp1479 = mem_1[tmp1447];
    assign tmp1624 = {const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0, const1623_0};
    assign tmp1308 = {tmp1307, tmp1211};
    assign tmp190 = {shifted_w31[16], shifted_w31[17], shifted_w31[18], shifted_w31[19], shifted_w31[20], shifted_w31[21], shifted_w31[22], shifted_w31[23]};
    assign temp_32 = new_9;
    assign tmp777 = {const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0, const776_0};
    assign concat_w23 = tmp153;
        assign tmp970 = mem_3[tmp916];
    assign tmp2341 = tmp2357;
        assign tmp1982 = mem_4[tmp1807];
    assign tmp1979 = tmp1975 ^ tmp1978;
    assign tmp1250 = {tmp1249[0], tmp1249[1], tmp1249[2], tmp1249[3], tmp1249[4], tmp1249[5], tmp1249[6], tmp1249[7]};
    assign tmp2070 = {temp_25[112], temp_25[113], temp_25[114], temp_25[115], temp_25[116], temp_25[117], temp_25[118], temp_25[119]};
        assign tmp1701 = mem_4[tmp1515];
    assign tmp266 = {new_state[88], new_state[89], new_state[90], new_state[91], new_state[92], new_state[93], new_state[94], new_state[95]};
    assign b3_w15 = tmp91;
    assign tmp160 = {tmp158[16], tmp158[17], tmp158[18], tmp158[19], tmp158[20], tmp158[21], tmp158[22], tmp158[23]};
    assign tmp470 = tmp468 ^ tmp469;
    assign tmp1727 = {temp_20[120], temp_20[121], temp_20[122], temp_20[123], temp_20[124], temp_20[125], temp_20[126], temp_20[127]};
    assign tmp943 = tmp1113;
    assign tmp1658 = tmp1654 ^ tmp1657;
    assign tmp91 = {shifted_w15[8], shifted_w15[9], shifted_w15[10], shifted_w15[11], shifted_w15[12], shifted_w15[13], shifted_w15[14], shifted_w15[15]};
    assign tmp178 = {rc1_w27, rc2_w27, rc3_w27, rc4_w27};
    assign tmp2165 = {tmp2164[0], tmp2164[1], tmp2164[2], tmp2164[3], tmp2164[4], tmp2164[5], tmp2164[6], tmp2164[7]};
    assign tmp1265 = tmp1263 ^ tmp1264;
        assign tmp1359 = mem_3[tmp1217];
    assign tmp2465 = tmp2461 ^ tmp2464;
        assign tmp306 = mem_1[tmp274];
    assign shifted_w11 = tmp63;
        assign tmp2647 = mem_1[tmp2615];
    assign rc2_w31 = const200_0;
    assign tmp2724 = {const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0, const2723_0};
    assign tmp1028 = tmp1024 ^ tmp1027;
    assign tmp6 = {aes_key[64], aes_key[65], aes_key[66], aes_key[67], aes_key[68], aes_key[69], aes_key[70], aes_key[71], aes_key[72], aes_key[73], aes_key[74], aes_key[75], aes_key[76], aes_key[77], aes_key[78], aes_key[79], aes_key[80], aes_key[81], aes_key[82], aes_key[83], aes_key[84], aes_key[85], aes_key[86], aes_key[87], aes_key[88], aes_key[89], aes_key[90], aes_key[91], aes_key[92], aes_key[93], aes_key[94], aes_key[95]};
    assign tmp347 = tmp407;
    assign new_state = new_1;
    assign tmp314 = {temp_1[96], temp_1[97], temp_1[98], temp_1[99], temp_1[100], temp_1[101], temp_1[102], temp_1[103]};
    assign tmp849 = {temp_8[112], temp_8[113], temp_8[114], temp_8[115], temp_8[116], temp_8[117], temp_8[118], temp_8[119]};
    assign concat_w39 = tmp253;
    assign tmp2634 = tmp2650;
    assign tmp2845 = {tmp2844, tmp2682};
    assign tmp2363 = {temp_29[112], temp_29[113], temp_29[114], temp_29[115], temp_29[116], temp_29[117], temp_29[118], temp_29[119]};
    assign tmp2410 = tmp2602;
    assign tmp2548 = {tmp2547, tmp2388};
    assign tmp419 = {tmp418[0], tmp418[1], tmp418[2], tmp418[3], tmp418[4], tmp418[5], tmp418[6], tmp418[7]};
    assign tmp2955 = {temp_37[64], temp_37[65], temp_37[66], temp_37[67], temp_37[68], temp_37[69], temp_37[70], temp_37[71]};
    assign tmp1527 = tmp1675;
    assign tmp611 = {temp_5[64], temp_5[65], temp_5[66], temp_5[67], temp_5[68], temp_5[69], temp_5[70], temp_5[71]};
    assign a2_w7 = tmp35;
    assign tmp951 = {tmp950, tmp916};
    assign tmp476 = {const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0, const475_0};
    assign tmp2116 = tmp2297;
    assign tmp2517 = tmp2513 ^ tmp2516;
    assign rc4_w35 = const227_0;
    assign tmp1436 = {temp_16[104], temp_16[105], temp_16[106], temp_16[107], temp_16[108], temp_16[109], temp_16[110], temp_16[111]};
    assign tmp2092 = {temp_26[72], temp_26[73], temp_26[74], temp_26[75], temp_26[76], temp_26[77], temp_26[78], temp_26[79]};
    assign tmp2146 = {const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0, const2145_0};
    assign tmp2196 = tmp2192 ^ tmp2195;
    assign tmp1804 = {temp_22[32], temp_22[33], temp_22[34], temp_22[35], temp_22[36], temp_22[37], temp_22[38], temp_22[39]};
    assign tmp1389 = tmp1385 ^ tmp1388;
    assign tmp571 = tmp587;
    assign tmp993 = {tmp992[0], tmp992[1], tmp992[2], tmp992[3], tmp992[4], tmp992[5], tmp992[6], tmp992[7]};
    assign new_1 = tmp261;
        assign tmp194 = mem_1[b2_w31];
    assign tmp2964 = {tmp2948, tmp2953, tmp2958, tmp2963, tmp2952, tmp2957, tmp2962, tmp2951, tmp2956, tmp2961, tmp2950, tmp2955, tmp2960, tmp2949, tmp2954, tmp2959};
    assign tmp497 = {tmp496, tmp337};
    assign tmp624 = {temp_6[96], temp_6[97], temp_6[98], temp_6[99], temp_6[100], temp_6[101], temp_6[102], temp_6[103]};
    assign tmp234 = {tmp233[24], tmp233[25], tmp233[26], tmp233[27], tmp233[28], tmp233[29], tmp233[30], tmp233[31]};
    assign tmp1235 = tmp1394;
    assign tmp1441 = {temp_16[64], temp_16[65], temp_16[66], temp_16[67], temp_16[68], temp_16[69], temp_16[70], temp_16[71]};
        assign tmp1761 = mem_1[tmp1729];
    assign tmp235 = {tmp233[16], tmp233[17], tmp233[18], tmp233[19], tmp233[20], tmp233[21], tmp233[22], tmp233[23]};
    assign tmp357 = tmp527;
        assign tmp119 = mem_1[b2_w19];
    assign tmp2385 = {temp_30[72], temp_30[73], temp_30[74], temp_30[75], temp_30[76], temp_30[77], temp_30[78], temp_30[79]};
    assign tmp1166 = tmp1182;
    assign tmp558 = {temp_4[96], temp_4[97], temp_4[98], temp_4[99], temp_4[100], temp_4[101], temp_4[102], temp_4[103]};
    assign tmp1462 = tmp1478;
    assign temp_29 = tmp2361;
    assign tmp2541 = tmp2537 ^ tmp2540;
    assign tmp453 = {tmp452, tmp334};
    assign a3_w15 = tmp86;
    assign tmp2455 = {const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0, const2454_0};
    assign tmp156 = tmp155 ^ tmp131;
    assign tmp1950 = {tmp1949, tmp1801};
    assign tmp2680 = {temp_34[56], temp_34[57], temp_34[58], temp_34[59], temp_34[60], temp_34[61], temp_34[62], temp_34[63]};
    assign tmp1890 = {tmp1889, tmp1800};
    assign tmp631 = {temp_6[40], temp_6[41], temp_6[42], temp_6[43], temp_6[44], temp_6[45], temp_6[46], temp_6[47]};
        assign tmp1640 = mem_3[tmp1509];
    assign tmp1612 = {const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0, const1611_0};
    assign tmp1830 = {tmp1829, tmp1795};
    assign tmp974 = {const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0, const973_0};
    assign tmp1824 = tmp2016;
        assign tmp1055 = mem_4[tmp924];
    assign tmp1954 = {tmp1953, tmp1802};
    assign tmp2329 = tmp2345;
    assign tmp2877 = {tmp2876, tmp2684};
    assign tmp1485 = {temp_17[104], temp_17[105], temp_17[106], temp_17[107], temp_17[108], temp_17[109], temp_17[110], temp_17[111]};
    assign tmp801 = {const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0, const800_0};
    assign tmp1059 = {tmp1058, tmp925};
    assign tmp2505 = tmp2501 ^ tmp2504;
    assign tmp2379 = {temp_30[120], temp_30[121], temp_30[122], temp_30[123], temp_30[124], temp_30[125], temp_30[126], temp_30[127]};
        assign tmp2412 = mem_4[tmp2380];
    assign tmp1992 = {tmp1991[0], tmp1991[1], tmp1991[2], tmp1991[3], tmp1991[4], tmp1991[5], tmp1991[6], tmp1991[7]};
    assign tmp1020 = tmp1018 ^ tmp1019;
    assign tmp1789 = {temp_21[16], temp_21[17], temp_21[18], temp_21[19], temp_21[20], temp_21[21], temp_21[22], temp_21[23]};
    assign tmp2559 = {const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0, const2558_0};
    assign tmp1634 = tmp1630 ^ tmp1633;
        assign tmp1090 = mem_3[tmp926];
    assign tmp1800 = {temp_22[64], temp_22[65], temp_22[66], temp_22[67], temp_22[68], temp_22[69], temp_22[70], temp_22[71]};
    assign tmp841 = {const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0, const840_0};
    assign tmp2710 = tmp2706 ^ tmp2709;
    assign tmp1552 = {const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0, const1551_0};
    assign xor_w7 = tmp54;
    assign tmp2023 = {temp_24[96], temp_24[97], temp_24[98], temp_24[99], temp_24[100], temp_24[101], temp_24[102], temp_24[103]};
    assign rc3_w27 = const176_0;
        assign tmp1849 = mem_3[tmp1795];
    assign tmp854 = {temp_8[72], temp_8[73], temp_8[74], temp_8[75], temp_8[76], temp_8[77], temp_8[78], temp_8[79]};
    assign tmp2236 = tmp2232 ^ tmp2235;
    assign tmp1416 = {tmp1415, tmp1220};
    assign tmp17 = {shifted_w3[0], shifted_w3[1], shifted_w3[2], shifted_w3[3], shifted_w3[4], shifted_w3[5], shifted_w3[6], shifted_w3[7]};
    assign b4_w23 = tmp142;
    assign tmp2392 = {temp_30[16], temp_30[17], temp_30[18], temp_30[19], temp_30[20], temp_30[21], temp_30[22], temp_30[23]};
    assign tmp1149 = {temp_12[56], temp_12[57], temp_12[58], temp_12[59], temp_12[60], temp_12[61], temp_12[62], temp_12[63]};
    assign tmp850 = {temp_8[104], temp_8[105], temp_8[106], temp_8[107], temp_8[108], temp_8[109], temp_8[110], temp_8[111]};
    assign tmp2675 = {temp_34[96], temp_34[97], temp_34[98], temp_34[99], temp_34[100], temp_34[101], temp_34[102], temp_34[103]};
        assign tmp1581 = mem_4[tmp1505];
    assign tmp1553 = {tmp1552, tmp1500};
    assign tmp1788 = {temp_21[24], temp_21[25], temp_21[26], temp_21[27], temp_21[28], temp_21[29], temp_21[30], temp_21[31]};
    assign substituted_w3 = tmp22;
        assign tmp2860 = mem_3[tmp2685];
    assign rc1_w23 = tmp149;
    assign tmp1487 = {temp_17[88], temp_17[89], temp_17[90], temp_17[91], temp_17[92], temp_17[93], temp_17[94], temp_17[95]};
    assign temp_14 = tmp1206;
    assign tmp2748 = {const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0, const2747_0};
    assign tmp633 = {temp_6[24], temp_6[25], temp_6[26], temp_6[27], temp_6[28], temp_6[29], temp_6[30], temp_6[31]};
    assign tmp1740 = {temp_20[16], temp_20[17], temp_20[18], temp_20[19], temp_20[20], temp_20[21], temp_20[22], temp_20[23]};
    assign tmp2637 = tmp2653;
    assign tmp2906 = {temp_36[64], temp_36[65], temp_36[66], temp_36[67], temp_36[68], temp_36[69], temp_36[70], temp_36[71]};
    assign tmp1334 = {tmp1333[0], tmp1333[1], tmp1333[2], tmp1333[3], tmp1333[4], tmp1333[5], tmp1333[6], tmp1333[7]};
    assign tmp1437 = {temp_16[96], temp_16[97], temp_16[98], temp_16[99], temp_16[100], temp_16[101], temp_16[102], temp_16[103]};
        assign tmp529 = mem_4[tmp343];
    assign tmp283 = tmp299;
    assign tmp2687 = {temp_34[0], temp_34[1], temp_34[2], temp_34[3], temp_34[4], temp_34[5], temp_34[6], temp_34[7]};
    assign tmp2904 = {temp_36[80], temp_36[81], temp_36[82], temp_36[83], temp_36[84], temp_36[85], temp_36[86], temp_36[87]};
    assign tmp209 = {tmp208[24], tmp208[25], tmp208[26], tmp208[27], tmp208[28], tmp208[29], tmp208[30], tmp208[31]};
    assign tmp2880 = {const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0, const2879_0};
    assign tmp53 = {rc1_w7, rc2_w7, rc3_w7, rc4_w7};
    assign tmp136 = {tmp133[8], tmp133[9], tmp133[10], tmp133[11], tmp133[12], tmp133[13], tmp133[14], tmp133[15]};
    assign tmp1872 = {tmp1871[0], tmp1871[1], tmp1871[2], tmp1871[3], tmp1871[4], tmp1871[5], tmp1871[6], tmp1871[7]};
        assign tmp2705 = mem_4[tmp2673];
    assign tmp1284 = {tmp1283, tmp1209};
    assign tmp2688 = tmp2715;
        assign tmp1628 = mem_3[tmp1508];
    assign tmp1247 = {const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0, const1246_0};
    assign temp_16 = new_5;
        assign tmp1556 = mem_3[tmp1502];
    assign tmp755 = tmp751 ^ tmp754;
    assign tmp2003 = tmp1999 ^ tmp2002;
    assign tmp1836 = {tmp1835[0], tmp1835[1], tmp1835[2], tmp1835[3], tmp1835[4], tmp1835[5], tmp1835[6], tmp1835[7]};
    assign b4_w31 = tmp192;
    assign tmp910 = {temp_9[16], temp_9[17], temp_9[18], temp_9[19], temp_9[20], temp_9[21], temp_9[22], temp_9[23]};
        assign tmp301 = mem_1[tmp269];
    assign tmp1012 = tmp1008 ^ tmp1011;
    assign tmp2321 = {temp_28[56], temp_28[57], temp_28[58], temp_28[59], temp_28[60], temp_28[61], temp_28[62], temp_28[63]};
    assign tmp1947 = tmp1945 ^ tmp1946;
    assign tmp464 = {const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0, const463_0};
    assign tmp2699 = tmp2847;
    assign tmp791 = tmp787 ^ tmp790;
    assign tmp779 = tmp775 ^ tmp778;
    assign tmp1508 = {temp_18[56], temp_18[57], temp_18[58], temp_18[59], temp_18[60], temp_18[61], temp_18[62], temp_18[63]};
    assign tmp65 = {shifted_w11[16], shifted_w11[17], shifted_w11[18], shifted_w11[19], shifted_w11[20], shifted_w11[21], shifted_w11[22], shifted_w11[23]};
    assign tmp2395 = tmp2422;
    assign tmp1215 = {temp_14[56], temp_14[57], temp_14[58], temp_14[59], temp_14[60], temp_14[61], temp_14[62], temp_14[63]};
        assign tmp299 = mem_1[tmp267];
        assign tmp1473 = mem_1[tmp1441];
    assign tmp1304 = {tmp1303, tmp1214};
    assign tmp2332 = tmp2348;
        assign tmp1324 = mem_4[tmp1211];
    assign tmp288 = tmp304;
    assign tmp1455 = tmp1471;
    assign tmp2456 = {tmp2455, tmp2381};
    assign tmp2150 = {const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0, const2149_0};
    assign tmp2853 = {tmp2852, tmp2686};
    assign tmp2342 = tmp2358;
    assign tmp615 = {temp_5[32], temp_5[33], temp_5[34], temp_5[35], temp_5[36], temp_5[37], temp_5[38], temp_5[39]};
        assign tmp49 = mem_2[const48_2];
    assign tmp2714 = tmp2710 ^ tmp2713;
    assign tmp813 = {const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0, const812_0};
    assign tmp2224 = tmp2220 ^ tmp2223;
    assign tmp1140 = temp_11 ^ tmp1139;
        assign tmp1287 = mem_3[tmp1211];
    assign tmp2615 = {temp_32[48], temp_32[49], temp_32[50], temp_32[51], temp_32[52], temp_32[53], temp_32[54], temp_32[55]};
    assign tmp1594 = tmp1592 ^ tmp1593;
    assign tmp2324 = {temp_28[32], temp_28[33], temp_28[34], temp_28[35], temp_28[36], temp_28[37], temp_28[38], temp_28[39]};
    assign tmp2745 = {tmp2744, tmp2673};
    assign tmp2918 = tmp2934;
    assign tmp2506 = {tmp2505[0], tmp2505[1], tmp2505[2], tmp2505[3], tmp2505[4], tmp2505[5], tmp2505[6], tmp2505[7]};
    assign tmp14 = {shifted_w3[24], shifted_w3[25], shifted_w3[26], shifted_w3[27], shifted_w3[28], shifted_w3[29], shifted_w3[30], shifted_w3[31]};
        assign tmp2351 = mem_1[tmp2319];
    assign a1_w31 = tmp184;
    assign tmp2083 = {temp_25[8], temp_25[9], temp_25[10], temp_25[11], temp_25[12], temp_25[13], temp_25[14], temp_25[15]};
    assign tmp607 = {temp_5[96], temp_5[97], temp_5[98], temp_5[99], temp_5[100], temp_5[101], temp_5[102], temp_5[103]};
    assign tmp2194 = {const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0, const2193_0};
    assign tmp2513 = tmp2509 ^ tmp2512;
    assign tmp280 = tmp296;
    assign w4 = tmp30;
    assign tmp381 = {tmp380, tmp328};
    assign tmp2431 = {const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0, const2430_0};
    assign tmp1244 = {tmp1243, tmp1209};
    assign tmp2372 = {temp_29[40], temp_29[41], temp_29[42], temp_29[43], temp_29[44], temp_29[45], temp_29[46], temp_29[47]};
    assign tmp333 = {temp_2[80], temp_2[81], temp_2[82], temp_2[83], temp_2[84], temp_2[85], temp_2[86], temp_2[87]};
    assign tmp1313 = tmp1311 ^ tmp1312;
    assign tmp1003 = {tmp1002, tmp921};
    assign tmp2485 = tmp2483 ^ tmp2484;
    assign tmp1572 = {const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0, const1571_0};
    assign tmp1164 = tmp1180;
    assign tmp1675 = {tmp1674[0], tmp1674[1], tmp1674[2], tmp1674[3], tmp1674[4], tmp1674[5], tmp1674[6], tmp1674[7]};
    assign tmp1218 = {temp_14[32], temp_14[33], temp_14[34], temp_14[35], temp_14[36], temp_14[37], temp_14[38], temp_14[39]};
    assign tmp2302 = {const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0, const2301_0};
    assign a2_w3 = tmp10;
    assign tmp991 = {tmp990, tmp916};
        assign tmp1641 = mem_4[tmp1510];
    assign input_wire_11 = temp_38;
    assign tmp2535 = {const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0, const2534_0};
    assign b3_w11 = tmp66;
    assign tmp2518 = {tmp2517[0], tmp2517[1], tmp2517[2], tmp2517[3], tmp2517[4], tmp2517[5], tmp2517[6], tmp2517[7]};
    assign tmp1494 = {temp_17[32], temp_17[33], temp_17[34], temp_17[35], temp_17[36], temp_17[37], temp_17[38], temp_17[39]};
    assign tmp1084 = tmp1080 ^ tmp1083;
    assign tmp358 = tmp539;
    assign tmp552 = {tmp344, tmp345, tmp346, tmp347, tmp348, tmp349, tmp350, tmp351, tmp352, tmp353, tmp354, tmp355, tmp356, tmp357, tmp358, tmp359};
    assign tmp1943 = tmp1939 ^ tmp1942;
    assign tmp2080 = {temp_25[32], temp_25[33], temp_25[34], temp_25[35], temp_25[36], temp_25[37], temp_25[38], temp_25[39]};
    assign tmp2725 = {tmp2724, tmp2672};
    assign tmp915 = {temp_10[112], temp_10[113], temp_10[114], temp_10[115], temp_10[116], temp_10[117], temp_10[118], temp_10[119]};
    assign tmp2597 = tmp2593 ^ tmp2596;
    assign tmp265 = {new_state[96], new_state[97], new_state[98], new_state[99], new_state[100], new_state[101], new_state[102], new_state[103]};
    assign tmp2842 = tmp2838 ^ tmp2841;
    assign tmp1505 = {temp_18[80], temp_18[81], temp_18[82], temp_18[83], temp_18[84], temp_18[85], temp_18[86], temp_18[87]};
    assign tmp1315 = {const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0, const1314_0};
    assign b4_w11 = tmp67;
    assign tmp1484 = {temp_17[112], temp_17[113], temp_17[114], temp_17[115], temp_17[116], temp_17[117], temp_17[118], temp_17[119]};
    assign temp_21 = tmp1775;
    assign tmp2552 = {tmp2551, tmp2389};
    assign tmp440 = {const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0, const439_0};
        assign tmp1945 = mem_3[tmp1803];
    assign tmp62 = {tmp58[0], tmp58[1], tmp58[2], tmp58[3], tmp58[4], tmp58[5], tmp58[6], tmp58[7]};
    assign tmp1573 = {tmp1572, tmp1501};
    assign tmp491 = {tmp490[0], tmp490[1], tmp490[2], tmp490[3], tmp490[4], tmp490[5], tmp490[6], tmp490[7]};
    assign tmp1204 = {temp_13[8], temp_13[9], temp_13[10], temp_13[11], temp_13[12], temp_13[13], temp_13[14], temp_13[15]};
    assign tmp1744 = tmp1760;
        assign tmp833 = mem_3[tmp636];
        assign tmp1019 = mem_4[tmp921];
    assign tmp873 = tmp889;
    assign tmp2034 = {temp_24[8], temp_24[9], temp_24[10], temp_24[11], temp_24[12], temp_24[13], temp_24[14], temp_24[15]};
    assign tmp1534 = tmp1532 ^ tmp1533;
    assign tmp1104 = tmp1102 ^ tmp1103;
        assign tmp774 = mem_4[tmp632];
        assign tmp2638 = mem_1[tmp2606];
        assign tmp594 = mem_1[tmp562];
    assign tmp1365 = tmp1361 ^ tmp1364;
    assign tmp1966 = {tmp1965, tmp1803};
        assign tmp1470 = mem_1[tmp1438];
    assign tmp643 = tmp736;
    assign tmp1267 = {const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0, const1266_0};
    assign tmp1579 = {tmp1578[0], tmp1578[1], tmp1578[2], tmp1578[3], tmp1578[4], tmp1578[5], tmp1578[6], tmp1578[7]};
        assign tmp2346 = mem_1[tmp2314];
        assign tmp1079 = mem_4[tmp922];
        assign tmp2836 = mem_3[tmp2683];
    assign tmp2001 = {const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0, const2000_0};
    assign tmp2545 = tmp2543 ^ tmp2544;
    assign tmp1205 = {temp_13[0], temp_13[1], temp_13[2], temp_13[3], temp_13[4], temp_13[5], temp_13[6], temp_13[7]};
        assign tmp2347 = mem_1[tmp2315];
    assign tmp667 = tmp665 ^ tmp666;
    assign tmp2090 = {temp_26[88], temp_26[89], temp_26[90], temp_26[91], temp_26[92], temp_26[93], temp_26[94], temp_26[95]};
    assign tmp1211 = {temp_14[88], temp_14[89], temp_14[90], temp_14[91], temp_14[92], temp_14[93], temp_14[94], temp_14[95]};
    assign tmp1794 = {temp_22[112], temp_22[113], temp_22[114], temp_22[115], temp_22[116], temp_22[117], temp_22[118], temp_22[119]};
    assign tmp1516 = tmp1543;
    assign rc2_w11 = const75_0;
    assign tmp63 = {a2_w11, a3_w11, a4_w11, a1_w11};
    assign c4_w11 = tmp71;
    assign tmp1370 = {tmp1369[0], tmp1369[1], tmp1369[2], tmp1369[3], tmp1369[4], tmp1369[5], tmp1369[6], tmp1369[7]};
    assign tmp584 = tmp600;
    assign tmp1369 = tmp1365 ^ tmp1368;
    assign tmp2564 = {tmp2563, tmp2394};
    assign tmp610 = {temp_5[72], temp_5[73], temp_5[74], temp_5[75], temp_5[76], temp_5[77], temp_5[78], temp_5[79]};
    assign tmp92 = {shifted_w15[0], shifted_w15[1], shifted_w15[2], shifted_w15[3], shifted_w15[4], shifted_w15[5], shifted_w15[6], shifted_w15[7]};
    assign tmp574 = tmp590;
        assign tmp884 = mem_1[tmp852];
    assign tmp1493 = {temp_17[40], temp_17[41], temp_17[42], temp_17[43], temp_17[44], temp_17[45], temp_17[46], temp_17[47]};
    assign tmp1086 = {const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0, const1085_0};
    assign tmp2826 = tmp2824 ^ tmp2825;
    assign tmp1273 = tmp1269 ^ tmp1272;
    assign tmp2440 = {tmp2439, tmp2379};
    assign tmp2189 = {tmp2188[0], tmp2188[1], tmp2188[2], tmp2188[3], tmp2188[4], tmp2188[5], tmp2188[6], tmp2188[7]};
    assign tmp2577 = tmp2573 ^ tmp2576;
    assign tmp1206 = {tmp1190, tmp1195, tmp1200, tmp1205, tmp1194, tmp1199, tmp1204, tmp1193, tmp1198, tmp1203, tmp1192, tmp1197, tmp1202, tmp1191, tmp1196, tmp1201};
    assign tmp2327 = {temp_28[8], temp_28[9], temp_28[10], temp_28[11], temp_28[12], temp_28[13], temp_28[14], temp_28[15]};
    assign tmp1597 = {tmp1596, tmp1507};
    assign tmp1120 = tmp1116 ^ tmp1119;
    assign tmp472 = {const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0, const471_0};
    assign tmp534 = tmp530 ^ tmp533;
    assign tmp159 = {tmp158[24], tmp158[25], tmp158[26], tmp158[27], tmp158[28], tmp158[29], tmp158[30], tmp158[31]};
    assign tmp685 = {const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0, const684_0};
    assign tmp2626 = tmp2642;
    assign tmp556 = {temp_4[112], temp_4[113], temp_4[114], temp_4[115], temp_4[116], temp_4[117], temp_4[118], temp_4[119]};
    assign tmp1452 = tmp1468;
    assign tmp1692 = {const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0, const1691_0};
        assign tmp1188 = mem_1[tmp1156];
        assign tmp2717 = mem_4[tmp2674];
    assign a1_w11 = tmp59;
    assign c3_w27 = tmp170;
        assign tmp121 = mem_1[b4_w19];
    assign c2_w7 = tmp44;
    assign tmp2376 = {temp_29[8], temp_29[9], temp_29[10], temp_29[11], temp_29[12], temp_29[13], temp_29[14], temp_29[15]};
    assign c3_w23 = tmp145;
    assign tmp878 = tmp894;
        assign tmp2848 = mem_3[tmp2684];
    assign tmp612 = {temp_5[56], temp_5[57], temp_5[58], temp_5[59], temp_5[60], temp_5[61], temp_5[62], temp_5[63]};
    assign tmp229 = concat_w35 ^ substituted_w35;
    assign tmp2553 = tmp2549 ^ tmp2552;
    assign tmp2446 = {tmp2445[0], tmp2445[1], tmp2445[2], tmp2445[3], tmp2445[4], tmp2445[5], tmp2445[6], tmp2445[7]};
    assign tmp2369 = {temp_29[64], temp_29[65], temp_29[66], temp_29[67], temp_29[68], temp_29[69], temp_29[70], temp_29[71]};
    assign tmp710 = {tmp709, tmp628};
    assign tmp2623 = tmp2639;
    assign tmp2607 = {temp_32[112], temp_32[113], temp_32[114], temp_32[115], temp_32[116], temp_32[117], temp_32[118], temp_32[119]};
    assign tmp1546 = tmp1544 ^ tmp1545;
    assign tmp185 = {tmp183[16], tmp183[17], tmp183[18], tmp183[19], tmp183[20], tmp183[21], tmp183[22], tmp183[23]};
    assign tmp142 = {shifted_w23[0], shifted_w23[1], shifted_w23[2], shifted_w23[3], shifted_w23[4], shifted_w23[5], shifted_w23[6], shifted_w23[7]};
    assign tmp1863 = tmp1861 ^ tmp1862;
    assign tmp2706 = tmp2704 ^ tmp2705;
    assign tmp1388 = {tmp1387, tmp1221};
    assign tmp2686 = {temp_34[8], temp_34[9], temp_34[10], temp_34[11], temp_34[12], temp_34[13], temp_34[14], temp_34[15]};
        assign tmp653 = mem_3[tmp621];
    assign tmp688 = {tmp687[0], tmp687[1], tmp687[2], tmp687[3], tmp687[4], tmp687[5], tmp687[6], tmp687[7]};
    assign tmp2282 = {const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0, const2281_0};
    assign tmp1878 = {tmp1877, tmp1799};
    assign tmp11 = {w3[8], w3[9], w3[10], w3[11], w3[12], w3[13], w3[14], w3[15]};
        assign tmp1007 = mem_4[tmp920];
    assign tmp963 = {tmp962, tmp917};
    assign a1_w39 = tmp234;
    assign tmp1074 = {const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0, const1073_0};
    assign tmp803 = tmp799 ^ tmp802;
    assign tmp2858 = tmp2854 ^ tmp2857;
    assign tmp832 = {tmp831[0], tmp831[1], tmp831[2], tmp831[3], tmp831[4], tmp831[5], tmp831[6], tmp831[7]};
    assign tmp2966 = temp_38 ^ tmp2965;
        assign tmp2190 = mem_3[tmp2092];
    assign tmp1891 = tmp1887 ^ tmp1890;
    assign tmp189 = {shifted_w31[24], shifted_w31[25], shifted_w31[26], shifted_w31[27], shifted_w31[28], shifted_w31[29], shifted_w31[30], shifted_w31[31]};
    assign tmp605 = {temp_5[112], temp_5[113], temp_5[114], temp_5[115], temp_5[116], temp_5[117], temp_5[118], temp_5[119]};
        assign tmp1474 = mem_1[tmp1442];
    assign tmp918 = {temp_10[88], temp_10[89], temp_10[90], temp_10[91], temp_10[92], temp_10[93], temp_10[94], temp_10[95]};
    assign tmp2397 = tmp2446;
    assign tmp1786 = {temp_21[40], temp_21[41], temp_21[42], temp_21[43], temp_21[44], temp_21[45], temp_21[46], temp_21[47]};
    assign tmp217 = {shifted_w35[0], shifted_w35[1], shifted_w35[2], shifted_w35[3], shifted_w35[4], shifted_w35[5], shifted_w35[6], shifted_w35[7]};
    assign tmp2576 = {tmp2575, tmp2391};
    assign tmp16 = {shifted_w3[8], shifted_w3[9], shifted_w3[10], shifted_w3[11], shifted_w3[12], shifted_w3[13], shifted_w3[14], shifted_w3[15]};
    assign tmp232 = tmp231 ^ tmp207;
    assign tmp2557 = tmp2555 ^ tmp2556;
    assign tmp748 = {tmp747[0], tmp747[1], tmp747[2], tmp747[3], tmp747[4], tmp747[5], tmp747[6], tmp747[7]};
        assign tmp1348 = mem_4[tmp1217];
    assign tmp1146 = {temp_12[80], temp_12[81], temp_12[82], temp_12[83], temp_12[84], temp_12[85], temp_12[86], temp_12[87]};
    assign tmp1035 = {tmp1034, tmp919};
    assign tmp2601 = tmp2597 ^ tmp2600;
        assign tmp2287 = mem_4[tmp2101];
    assign tmp2014 = {tmp2013, tmp1807};
    assign a4_w19 = tmp112;
    assign substituted_w7 = tmp47;
    assign tmp1548 = {const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0, const1547_0};
    assign tmp2427 = {const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0, const2426_0};
    assign tmp874 = tmp890;
    assign tmp563 = {temp_4[56], temp_4[57], temp_4[58], temp_4[59], temp_4[60], temp_4[61], temp_4[62], temp_4[63]};
    assign tmp1128 = tmp1126 ^ tmp1127;
    assign tmp2829 = {tmp2828, tmp2680};
        assign tmp880 = mem_1[tmp848];
    assign tmp1000 = tmp996 ^ tmp999;
    assign tmp1601 = {tmp1600, tmp1504};
    assign tmp2797 = {tmp2796, tmp2678};
    assign tmp1460 = tmp1476;
    assign tmp2389 = {temp_30[40], temp_30[41], temp_30[42], temp_30[43], temp_30[44], temp_30[45], temp_30[46], temp_30[47]};
    assign tmp2578 = {tmp2577[0], tmp2577[1], tmp2577[2], tmp2577[3], tmp2577[4], tmp2577[5], tmp2577[6], tmp2577[7]};
        assign tmp2424 = mem_4[tmp2381];
        assign tmp2202 = mem_3[tmp2093];
    assign tmp274 = {new_state[24], new_state[25], new_state[26], new_state[27], new_state[28], new_state[29], new_state[30], new_state[31]};
    assign tmp2106 = tmp2177;
    assign tmp2375 = {temp_29[16], temp_29[17], temp_29[18], temp_29[19], temp_29[20], temp_29[21], temp_29[22], temp_29[23]};
    assign tmp320 = {temp_1[48], temp_1[49], temp_1[50], temp_1[51], temp_1[52], temp_1[53], temp_1[54], temp_1[55]};
    assign b2_w35 = tmp215;
    assign tmp1062 = {const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0, const1061_0};
    assign tmp2038 = tmp2054;
    assign tmp2494 = {tmp2493[0], tmp2493[1], tmp2493[2], tmp2493[3], tmp2493[4], tmp2493[5], tmp2493[6], tmp2493[7]};
    assign tmp263 = {new_state[112], new_state[113], new_state[114], new_state[115], new_state[116], new_state[117], new_state[118], new_state[119]};
    assign tmp2662 = {temp_33[64], temp_33[65], temp_33[66], temp_33[67], temp_33[68], temp_33[69], temp_33[70], temp_33[71]};
    assign tmp606 = {temp_5[104], temp_5[105], temp_5[106], temp_5[107], temp_5[108], temp_5[109], temp_5[110], temp_5[111]};
        assign tmp2568 = mem_4[tmp2393];
    assign rc4_w3 = const27_0;
        assign tmp1126 = mem_3[tmp929];
        assign tmp308 = mem_1[tmp276];
    assign tmp2344 = tmp2360;
    assign tmp1320 = {tmp1319, tmp1212};
    assign tmp1687 = {tmp1686[0], tmp1686[1], tmp1686[2], tmp1686[3], tmp1686[4], tmp1686[5], tmp1686[6], tmp1686[7]};
    assign tmp345 = tmp383;
    assign tmp2682 = {temp_34[40], temp_34[41], temp_34[42], temp_34[43], temp_34[44], temp_34[45], temp_34[46], temp_34[47]};
    assign tmp819 = tmp815 ^ tmp818;
        assign tmp24 = mem_2[const23_1];
    assign tmp109 = {tmp108[24], tmp108[25], tmp108[26], tmp108[27], tmp108[28], tmp108[29], tmp108[30], tmp108[31]};
    assign temp_34 = tmp2671;
    assign tmp315 = {temp_1[88], temp_1[89], temp_1[90], temp_1[91], temp_1[92], temp_1[93], temp_1[94], temp_1[95]};
        assign tmp1408 = mem_4[tmp1222];
    assign tmp712 = {tmp711[0], tmp711[1], tmp711[2], tmp711[3], tmp711[4], tmp711[5], tmp711[6], tmp711[7]};
    assign tmp1831 = tmp1827 ^ tmp1830;
        assign tmp304 = mem_1[tmp272];
    assign tmp2312 = temp_27 ^ tmp2311;
        assign tmp1336 = mem_4[tmp1216];
        assign tmp2543 = mem_3[tmp2390];
    assign tmp905 = {temp_9[56], temp_9[57], temp_9[58], temp_9[59], temp_9[60], temp_9[61], temp_9[62], temp_9[63]};
    assign tmp1319 = {const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0, const1318_0};
        assign tmp2060 = mem_1[tmp2028];
    assign tmp2509 = tmp2507 ^ tmp2508;
    assign tmp1063 = {tmp1062, tmp922};
    assign tmp981 = {tmp980[0], tmp980[1], tmp980[2], tmp980[3], tmp980[4], tmp980[5], tmp980[6], tmp980[7]};
    assign tmp2480 = {tmp2479, tmp2383};
    assign tmp1072 = tmp1068 ^ tmp1071;
    assign tmp2228 = tmp2226 ^ tmp2227;
    assign tmp998 = {const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0, const997_0};
    assign tmp130 = tmp105 ^ xor_w19;
    assign tmp2852 = {const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0, const2851_0};
    assign tmp1316 = {tmp1315, tmp1211};
    assign temp_20 = new_6;
    assign c4_w39 = tmp246;
    assign tmp1023 = {tmp1022, tmp918};
    assign tmp1582 = tmp1580 ^ tmp1581;
    assign input_wire_7 = temp_23;
    assign tmp2016 = {tmp2015[0], tmp2015[1], tmp2015[2], tmp2015[3], tmp2015[4], tmp2015[5], tmp2015[6], tmp2015[7]};
    assign tmp57 = tmp56 ^ w6;
    assign rc3_w39 = const251_0;
    assign tmp1123 = {tmp1122, tmp927};
    assign tmp1364 = {tmp1363, tmp1215};
    assign tmp2266 = {const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0, const2265_0};
    assign b1_w31 = tmp189;
    assign tmp2669 = {temp_33[8], temp_33[9], temp_33[10], temp_33[11], temp_33[12], temp_33[13], temp_33[14], temp_33[15]};
        assign tmp193 = mem_1[b1_w31];
    assign tmp313 = {temp_1[104], temp_1[105], temp_1[106], temp_1[107], temp_1[108], temp_1[109], temp_1[110], temp_1[111]};
    assign tmp2962 = {temp_37[8], temp_37[9], temp_37[10], temp_37[11], temp_37[12], temp_37[13], temp_37[14], temp_37[15]};
        assign tmp2837 = mem_4[tmp2680];
    assign tmp542 = tmp540 ^ tmp541;
    assign tmp2670 = {temp_33[0], temp_33[1], temp_33[2], temp_33[3], temp_33[4], temp_33[5], temp_33[6], temp_33[7]};
    assign tmp1163 = tmp1179;
    assign tmp58 = tmp57 ^ w7;
    assign tmp2279 = {tmp2278, tmp2101};
    assign tmp1523 = tmp1627;
    assign tmp2156 = tmp2154 ^ tmp2155;
    assign tmp2199 = {tmp2198, tmp2091};
    assign tmp1609 = {tmp1608, tmp1504};
    assign tmp565 = {temp_4[40], temp_4[41], temp_4[42], temp_4[43], temp_4[44], temp_4[45], temp_4[46], temp_4[47]};
    assign tmp2108 = tmp2201;
    assign tmp1202 = {temp_13[24], temp_13[25], temp_13[26], temp_13[27], temp_13[28], temp_13[29], temp_13[30], temp_13[31]};
    assign tmp206 = tmp205 ^ tmp181;
    assign tmp814 = {tmp813, tmp636};
    assign tmp1440 = {temp_16[72], temp_16[73], temp_16[74], temp_16[75], temp_16[76], temp_16[77], temp_16[78], temp_16[79]};
    assign tmp1353 = tmp1349 ^ tmp1352;
    assign tmp1879 = tmp1875 ^ tmp1878;
    assign tmp1259 = {const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0, const1258_0};
    assign tmp1380 = {tmp1379, tmp1217};
    assign tmp2922 = tmp2938;
    assign tmp2888 = {const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0, const2887_0};
    assign tmp767 = tmp763 ^ tmp766;
        assign tmp468 = mem_3[tmp337];
    assign tmp1291 = {const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0, const1290_0};
    assign tmp59 = {tmp58[24], tmp58[25], tmp58[26], tmp58[27], tmp58[28], tmp58[29], tmp58[30], tmp58[31]};
    assign tmp1751 = tmp1767;
    assign c1_w31 = tmp193;
        assign tmp885 = mem_1[tmp853];
    assign tmp2309 = {tmp2308[0], tmp2308[1], tmp2308[2], tmp2308[3], tmp2308[4], tmp2308[5], tmp2308[6], tmp2308[7]};
        assign tmp2155 = mem_4[tmp2086];
        assign tmp1532 = mem_3[tmp1500];
    assign tmp2482 = {tmp2481[0], tmp2481[1], tmp2481[2], tmp2481[3], tmp2481[4], tmp2481[5], tmp2481[6], tmp2481[7]};
    assign tmp2632 = tmp2648;
    assign tmp1725 = {expanded_key[640], expanded_key[641], expanded_key[642], expanded_key[643], expanded_key[644], expanded_key[645], expanded_key[646], expanded_key[647], expanded_key[648], expanded_key[649], expanded_key[650], expanded_key[651], expanded_key[652], expanded_key[653], expanded_key[654], expanded_key[655], expanded_key[656], expanded_key[657], expanded_key[658], expanded_key[659], expanded_key[660], expanded_key[661], expanded_key[662], expanded_key[663], expanded_key[664], expanded_key[665], expanded_key[666], expanded_key[667], expanded_key[668], expanded_key[669], expanded_key[670], expanded_key[671], expanded_key[672], expanded_key[673], expanded_key[674], expanded_key[675], expanded_key[676], expanded_key[677], expanded_key[678], expanded_key[679], expanded_key[680], expanded_key[681], expanded_key[682], expanded_key[683], expanded_key[684], expanded_key[685], expanded_key[686], expanded_key[687], expanded_key[688], expanded_key[689], expanded_key[690], expanded_key[691], expanded_key[692], expanded_key[693], expanded_key[694], expanded_key[695], expanded_key[696], expanded_key[697], expanded_key[698], expanded_key[699], expanded_key[700], expanded_key[701], expanded_key[702], expanded_key[703], expanded_key[704], expanded_key[705], expanded_key[706], expanded_key[707], expanded_key[708], expanded_key[709], expanded_key[710], expanded_key[711], expanded_key[712], expanded_key[713], expanded_key[714], expanded_key[715], expanded_key[716], expanded_key[717], expanded_key[718], expanded_key[719], expanded_key[720], expanded_key[721], expanded_key[722], expanded_key[723], expanded_key[724], expanded_key[725], expanded_key[726], expanded_key[727], expanded_key[728], expanded_key[729], expanded_key[730], expanded_key[731], expanded_key[732], expanded_key[733], expanded_key[734], expanded_key[735], expanded_key[736], expanded_key[737], expanded_key[738], expanded_key[739], expanded_key[740], expanded_key[741], expanded_key[742], expanded_key[743], expanded_key[744], expanded_key[745], expanded_key[746], expanded_key[747], expanded_key[748], expanded_key[749], expanded_key[750], expanded_key[751], expanded_key[752], expanded_key[753], expanded_key[754], expanded_key[755], expanded_key[756], expanded_key[757], expanded_key[758], expanded_key[759], expanded_key[760], expanded_key[761], expanded_key[762], expanded_key[763], expanded_key[764], expanded_key[765], expanded_key[766], expanded_key[767]};
    assign tmp509 = {tmp508, tmp342};
    assign tmp1004 = tmp1000 ^ tmp1003;
    assign tmp2958 = {temp_37[40], temp_37[41], temp_37[42], temp_37[43], temp_37[44], temp_37[45], temp_37[46], temp_37[47]};
    assign temp_15 = tmp1431;
    assign tmp222 = {c1_w35, c2_w35, c3_w35, c4_w35};
    assign tmp731 = tmp727 ^ tmp730;
    assign tmp2841 = {tmp2840, tmp2681};
    assign tmp1101 = {tmp1100[0], tmp1100[1], tmp1100[2], tmp1100[3], tmp1100[4], tmp1100[5], tmp1100[6], tmp1100[7]};
    assign tmp2761 = {tmp2760, tmp2679};
    assign tmp1684 = {const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0, const1683_0};
    assign tmp721 = {const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0, const720_0};
    assign tmp2304 = tmp2300 ^ tmp2303;
    assign tmp2611 = {temp_32[80], temp_32[81], temp_32[82], temp_32[83], temp_32[84], temp_32[85], temp_32[86], temp_32[87]};
    assign tmp2322 = {temp_28[48], temp_28[49], temp_28[50], temp_28[51], temp_28[52], temp_28[53], temp_28[54], temp_28[55]};
    assign tmp365 = {tmp364, tmp330};
    assign tmp1884 = {tmp1883[0], tmp1883[1], tmp1883[2], tmp1883[3], tmp1883[4], tmp1883[5], tmp1883[6], tmp1883[7]};
    assign tmp55 = w4 ^ xor_w7;
    assign tmp1590 = tmp1586 ^ tmp1589;
    assign tmp1233 = tmp1370;
    assign tmp271 = {new_state[48], new_state[49], new_state[50], new_state[51], new_state[52], new_state[53], new_state[54], new_state[55]};
    assign tmp2044 = tmp2060;
    assign tmp2529 = tmp2525 ^ tmp2528;
    assign tmp1089 = {tmp1088[0], tmp1088[1], tmp1088[2], tmp1088[3], tmp1088[4], tmp1088[5], tmp1088[6], tmp1088[7]};
    assign tmp2738 = tmp2734 ^ tmp2737;
    assign tmp1622 = tmp1618 ^ tmp1621;
    assign c1_w39 = tmp243;
    assign tmp2949 = {temp_37[112], temp_37[113], temp_37[114], temp_37[115], temp_37[116], temp_37[117], temp_37[118], temp_37[119]};
    assign tmp341 = {temp_2[16], temp_2[17], temp_2[18], temp_2[19], temp_2[20], temp_2[21], temp_2[22], temp_2[23]};
    assign c3_w15 = tmp95;
    assign tmp329 = {temp_2[112], temp_2[113], temp_2[114], temp_2[115], temp_2[116], temp_2[117], temp_2[118], temp_2[119]};
    assign tmp1743 = tmp1759;
    assign tmp1639 = {tmp1638[0], tmp1638[1], tmp1638[2], tmp1638[3], tmp1638[4], tmp1638[5], tmp1638[6], tmp1638[7]};
    assign rc4_w23 = const152_0;
    assign tmp1405 = tmp1401 ^ tmp1404;
        assign tmp2058 = mem_1[tmp2026];
    assign tmp1295 = {const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0, const1294_0};
    assign c2_w23 = tmp144;
    assign tmp273 = {new_state[32], new_state[33], new_state[34], new_state[35], new_state[36], new_state[37], new_state[38], new_state[39]};
    assign tmp759 = tmp755 ^ tmp758;
    assign tmp275 = {new_state[16], new_state[17], new_state[18], new_state[19], new_state[20], new_state[21], new_state[22], new_state[23]};
        assign tmp1922 = mem_4[tmp1802];
    assign tmp2475 = {const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0, const2474_0};
    assign a3_w27 = tmp161;
    assign tmp1894 = {tmp1893, tmp1797};
    assign tmp846 = {expanded_key[1024], expanded_key[1025], expanded_key[1026], expanded_key[1027], expanded_key[1028], expanded_key[1029], expanded_key[1030], expanded_key[1031], expanded_key[1032], expanded_key[1033], expanded_key[1034], expanded_key[1035], expanded_key[1036], expanded_key[1037], expanded_key[1038], expanded_key[1039], expanded_key[1040], expanded_key[1041], expanded_key[1042], expanded_key[1043], expanded_key[1044], expanded_key[1045], expanded_key[1046], expanded_key[1047], expanded_key[1048], expanded_key[1049], expanded_key[1050], expanded_key[1051], expanded_key[1052], expanded_key[1053], expanded_key[1054], expanded_key[1055], expanded_key[1056], expanded_key[1057], expanded_key[1058], expanded_key[1059], expanded_key[1060], expanded_key[1061], expanded_key[1062], expanded_key[1063], expanded_key[1064], expanded_key[1065], expanded_key[1066], expanded_key[1067], expanded_key[1068], expanded_key[1069], expanded_key[1070], expanded_key[1071], expanded_key[1072], expanded_key[1073], expanded_key[1074], expanded_key[1075], expanded_key[1076], expanded_key[1077], expanded_key[1078], expanded_key[1079], expanded_key[1080], expanded_key[1081], expanded_key[1082], expanded_key[1083], expanded_key[1084], expanded_key[1085], expanded_key[1086], expanded_key[1087], expanded_key[1088], expanded_key[1089], expanded_key[1090], expanded_key[1091], expanded_key[1092], expanded_key[1093], expanded_key[1094], expanded_key[1095], expanded_key[1096], expanded_key[1097], expanded_key[1098], expanded_key[1099], expanded_key[1100], expanded_key[1101], expanded_key[1102], expanded_key[1103], expanded_key[1104], expanded_key[1105], expanded_key[1106], expanded_key[1107], expanded_key[1108], expanded_key[1109], expanded_key[1110], expanded_key[1111], expanded_key[1112], expanded_key[1113], expanded_key[1114], expanded_key[1115], expanded_key[1116], expanded_key[1117], expanded_key[1118], expanded_key[1119], expanded_key[1120], expanded_key[1121], expanded_key[1122], expanded_key[1123], expanded_key[1124], expanded_key[1125], expanded_key[1126], expanded_key[1127], expanded_key[1128], expanded_key[1129], expanded_key[1130], expanded_key[1131], expanded_key[1132], expanded_key[1133], expanded_key[1134], expanded_key[1135], expanded_key[1136], expanded_key[1137], expanded_key[1138], expanded_key[1139], expanded_key[1140], expanded_key[1141], expanded_key[1142], expanded_key[1143], expanded_key[1144], expanded_key[1145], expanded_key[1146], expanded_key[1147], expanded_key[1148], expanded_key[1149], expanded_key[1150], expanded_key[1151]};
    assign c4_w19 = tmp121;
    assign tmp1959 = tmp1957 ^ tmp1958;
    assign tmp1906 = {tmp1905, tmp1798};
    assign tmp1064 = tmp1060 ^ tmp1063;
    assign tmp2303 = {tmp2302, tmp2099};
    assign c2_w15 = tmp94;
    assign tmp386 = tmp384 ^ tmp385;
    assign tmp2089 = {temp_26[96], temp_26[97], temp_26[98], temp_26[99], temp_26[100], temp_26[101], temp_26[102], temp_26[103]};
        assign tmp1885 = mem_3[tmp1798];
    assign tmp2886 = tmp2884 ^ tmp2885;
    assign tmp172 = {c1_w27, c2_w27, c3_w27, c4_w27};
    assign tmp2832 = {const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0, const2831_0};
        assign tmp2054 = mem_1[tmp2022];
    assign tmp1080 = tmp1078 ^ tmp1079;
        assign tmp1688 = mem_3[tmp1513];
    assign tmp957 = {tmp956[0], tmp956[1], tmp956[2], tmp956[3], tmp956[4], tmp956[5], tmp956[6], tmp956[7]};
    assign tmp933 = tmp993;
    assign tmp770 = {tmp769, tmp629};
    assign tmp626 = {temp_6[80], temp_6[81], temp_6[82], temp_6[83], temp_6[84], temp_6[85], temp_6[86], temp_6[87]};
    assign substituted_w39 = tmp247;
    assign tmp2773 = {tmp2772, tmp2676};
    assign tmp2168 = tmp2166 ^ tmp2167;
    assign tmp1107 = {tmp1106, tmp929};
    assign tmp629 = {temp_6[56], temp_6[57], temp_6[58], temp_6[59], temp_6[60], temp_6[61], temp_6[62], temp_6[63]};
        assign tmp307 = mem_1[tmp275];
        assign tmp2057 = mem_1[tmp2025];
        assign tmp1593 = mem_4[tmp1506];
        assign tmp2448 = mem_4[tmp2379];
    assign tmp2170 = {const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0, const2169_0};
    assign tmp2296 = tmp2292 ^ tmp2295;
        assign tmp677 = mem_3[tmp623];
    assign tmp1636 = {const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0, const1635_0};
    assign tmp2328 = {temp_28[0], temp_28[1], temp_28[2], temp_28[3], temp_28[4], temp_28[5], temp_28[6], temp_28[7]};
    assign rc1_w3 = tmp24;
    assign tmp2381 = {temp_30[104], temp_30[105], temp_30[106], temp_30[107], temp_30[108], temp_30[109], temp_30[110], temp_30[111]};
    assign tmp81 = tmp80 ^ tmp56;
    assign tmp2449 = tmp2447 ^ tmp2448;
    assign tmp1498 = {temp_17[0], temp_17[1], temp_17[2], temp_17[3], temp_17[4], temp_17[5], temp_17[6], temp_17[7]};
    assign tmp1048 = tmp1044 ^ tmp1047;
    assign concat_w31 = tmp203;
    assign tmp1412 = {tmp1411, tmp1219};
    assign tmp1752 = tmp1768;
        assign tmp2357 = mem_1[tmp2325];
    assign tmp2628 = tmp2644;
    assign tmp2951 = {temp_37[96], temp_37[97], temp_37[98], temp_37[99], temp_37[100], temp_37[101], temp_37[102], temp_37[103]};
    assign tmp1919 = tmp1915 ^ tmp1918;
    assign tmp1194 = {temp_13[88], temp_13[89], temp_13[90], temp_13[91], temp_13[92], temp_13[93], temp_13[94], temp_13[95]};
    assign b4_w35 = tmp217;
    assign tmp945 = tmp1137;
    assign tmp137 = {tmp133[0], tmp133[1], tmp133[2], tmp133[3], tmp133[4], tmp133[5], tmp133[6], tmp133[7]};
    assign temp_9 = tmp896;
    assign tmp642 = tmp724;
    assign tmp1630 = tmp1628 ^ tmp1629;
    assign tmp1355 = {const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0, const1354_0};
        assign tmp1898 = mem_4[tmp1800];
        assign tmp360 = mem_3[tmp328];
        assign tmp761 = mem_3[tmp630];
    assign tmp823 = tmp821 ^ tmp822;
    assign tmp825 = {const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0, const824_0};
        assign tmp1420 = mem_4[tmp1219];
        assign tmp43 = mem_1[b1_w7];
    assign tmp404 = {const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0, const403_0};
    assign tmp2927 = tmp2943;
    assign tmp369 = {tmp368, tmp331};
    assign tmp586 = tmp602;
    assign tmp861 = {temp_8[16], temp_8[17], temp_8[18], temp_8[19], temp_8[20], temp_8[21], temp_8[22], temp_8[23]};
    assign tmp2331 = tmp2347;
    assign tmp1070 = {const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0, const1069_0};
    assign new_7 = tmp2019;
    assign tmp258 = tmp257 ^ tmp233;
    assign tmp521 = {tmp520, tmp343};
    assign tmp1584 = {const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0, const1583_0};
    assign tmp2659 = {temp_33[88], temp_33[89], temp_33[90], temp_33[91], temp_33[92], temp_33[93], temp_33[94], temp_33[95]};
    assign b3_w23 = tmp141;
    assign tmp1339 = {const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0, const1338_0};
        assign tmp1127 = mem_4[tmp926];
    assign tmp1784 = {temp_21[56], temp_21[57], temp_21[58], temp_21[59], temp_21[60], temp_21[61], temp_21[62], temp_21[63]};
    assign tmp1171 = tmp1187;
    assign tmp1491 = {temp_17[56], temp_17[57], temp_17[58], temp_17[59], temp_17[60], temp_17[61], temp_17[62], temp_17[63]};
    assign tmp1907 = tmp1903 ^ tmp1906;
    assign tmp2928 = tmp2944;
    assign tmp1618 = tmp1616 ^ tmp1617;
    assign tmp290 = tmp306;
    assign tmp1268 = {tmp1267, tmp1207};
    assign tmp484 = {const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0, const483_0};
    assign b2_w19 = tmp115;
        assign tmp1616 = mem_3[tmp1507];
    assign tmp2820 = {const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0, const2819_0};
    assign tmp374 = tmp372 ^ tmp373;
        assign tmp481 = mem_4[tmp339];
        assign tmp886 = mem_1[tmp854];
    assign tmp671 = tmp667 ^ tmp670;
    assign tmp2164 = tmp2160 ^ tmp2163;
        assign tmp2644 = mem_1[tmp2612];
    assign tmp2268 = tmp2264 ^ tmp2267;
    assign tmp104 = concat_w15 ^ substituted_w15;
    assign tmp1394 = {tmp1393[0], tmp1393[1], tmp1393[2], tmp1393[3], tmp1393[4], tmp1393[5], tmp1393[6], tmp1393[7]};
        assign tmp2639 = mem_1[tmp2607];
        assign tmp1174 = mem_1[tmp1142];
    assign tmp1736 = {temp_20[48], temp_20[49], temp_20[50], temp_20[51], temp_20[52], temp_20[53], temp_20[54], temp_20[55]};
    assign tmp2394 = {temp_30[0], temp_30[1], temp_30[2], temp_30[3], temp_30[4], temp_30[5], temp_30[6], temp_30[7]};
        assign tmp881 = mem_1[tmp849];
    assign tmp583 = tmp599;
    assign tmp1662 = tmp1658 ^ tmp1661;
    assign tmp2393 = {temp_30[8], temp_30[9], temp_30[10], temp_30[11], temp_30[12], temp_30[13], temp_30[14], temp_30[15]};
    assign tmp2285 = {tmp2284[0], tmp2284[1], tmp2284[2], tmp2284[3], tmp2284[4], tmp2284[5], tmp2284[6], tmp2284[7]};
    assign tmp2408 = tmp2578;
    assign tmp863 = {temp_8[0], temp_8[1], temp_8[2], temp_8[3], temp_8[4], temp_8[5], temp_8[6], temp_8[7]};
    assign tmp1379 = {const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0, const1378_0};
    assign rc3_w23 = const151_0;
    assign tmp705 = {const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0, const704_0};
    assign tmp2043 = tmp2059;
    assign tmp2585 = tmp2581 ^ tmp2584;
    assign tmp1731 = {temp_20[88], temp_20[89], temp_20[90], temp_20[91], temp_20[92], temp_20[93], temp_20[94], temp_20[95]};
    assign tmp2163 = {tmp2162, tmp2088};
    assign tmp2661 = {temp_33[72], temp_33[73], temp_33[74], temp_33[75], temp_33[76], temp_33[77], temp_33[78], temp_33[79]};
    assign tmp494 = tmp492 ^ tmp493;
    assign tmp862 = {temp_8[8], temp_8[9], temp_8[10], temp_8[11], temp_8[12], temp_8[13], temp_8[14], temp_8[15]};
    assign tmp2011 = tmp2007 ^ tmp2010;
        assign tmp2064 = mem_1[tmp2032];
    assign tmp1722 = tmp1718 ^ tmp1721;
    assign tmp673 = {const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0, const672_0};
    assign tmp1814 = tmp1896;
    assign tmp2715 = {tmp2714[0], tmp2714[1], tmp2714[2], tmp2714[3], tmp2714[4], tmp2714[5], tmp2714[6], tmp2714[7]};
        assign tmp1946 = mem_4[tmp1804];
    assign tmp327 = {tmp311, tmp316, tmp321, tmp326, tmp315, tmp320, tmp325, tmp314, tmp319, tmp324, tmp313, tmp318, tmp323, tmp312, tmp317, tmp322};
    assign b2_w23 = tmp140;
    assign tmp2763 = {tmp2762[0], tmp2762[1], tmp2762[2], tmp2762[3], tmp2762[4], tmp2762[5], tmp2762[6], tmp2762[7]};
    assign tmp1138 = {tmp930, tmp931, tmp932, tmp933, tmp934, tmp935, tmp936, tmp937, tmp938, tmp939, tmp940, tmp941, tmp942, tmp943, tmp944, tmp945};
    assign rc3_w15 = const101_0;
    assign tmp2195 = {tmp2194, tmp2090};
    assign tmp909 = {temp_9[24], temp_9[25], temp_9[26], temp_9[27], temp_9[28], temp_9[29], temp_9[30], temp_9[31]};
    assign tmp2524 = {tmp2523, tmp2390};
        assign tmp596 = mem_1[tmp564];
        assign tmp785 = mem_3[tmp632];
    assign tmp1213 = {temp_14[72], temp_14[73], temp_14[74], temp_14[75], temp_14[76], temp_14[77], temp_14[78], temp_14[79]};
    assign tmp1670 = tmp1666 ^ tmp1669;
    assign tmp1720 = {const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0, const1719_0};
    assign temp_33 = tmp2654;
    assign tmp1274 = {tmp1273[0], tmp1273[1], tmp1273[2], tmp1273[3], tmp1273[4], tmp1273[5], tmp1273[6], tmp1273[7]};
        assign tmp1677 = mem_4[tmp1513];
    assign tmp1356 = {tmp1355, tmp1215};
    assign tmp1729 = {temp_20[104], temp_20[105], temp_20[106], temp_20[107], temp_20[108], temp_20[109], temp_20[110], temp_20[111]};
    assign tmp436 = {const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0, const435_0};
    assign temp_8 = new_3;
    assign tmp843 = tmp839 ^ tmp842;
    assign tmp376 = {const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0, const375_0};
    assign substituted_w27 = tmp172;
        assign tmp2274 = mem_3[tmp2099];
    assign tmp811 = tmp809 ^ tmp810;
        assign tmp1993 = mem_3[tmp1807];
        assign tmp2286 = mem_3[tmp2100];
        assign tmp2131 = mem_4[tmp2088];
    assign tmp1506 = {temp_18[72], temp_18[73], temp_18[74], temp_18[75], temp_18[76], temp_18[77], temp_18[78], temp_18[79]};
    assign tmp1417 = tmp1413 ^ tmp1416;
    assign tmp164 = {shifted_w27[24], shifted_w27[25], shifted_w27[26], shifted_w27[27], shifted_w27[28], shifted_w27[29], shifted_w27[30], shifted_w27[31]};
    assign tmp1404 = {tmp1403, tmp1219};
        assign tmp245 = mem_1[b3_w39];
    assign rc2_w23 = const150_0;
        assign tmp1275 = mem_3[tmp1210];
    assign tmp807 = tmp803 ^ tmp806;
    assign temp_11 = tmp1138;
    assign tmp2794 = tmp2790 ^ tmp2793;
        assign tmp2250 = mem_3[tmp2097];
    assign tmp2869 = {tmp2868, tmp2684};
    assign tmp54 = concat_w7 ^ substituted_w7;
    assign tmp2013 = {const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0, const2012_0};
        assign tmp540 = mem_3[tmp343];
    assign tmp579 = tmp595;
    assign tmp1985 = {const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0, const1984_0};
    assign tmp418 = tmp414 ^ tmp417;
    assign tmp1051 = {tmp1050, tmp925};
    assign tmp2370 = {temp_29[56], temp_29[57], temp_29[58], temp_29[59], temp_29[60], temp_29[61], temp_29[62], temp_29[63]};
    assign tmp2921 = tmp2937;
    assign tmp2272 = tmp2268 ^ tmp2271;
        assign tmp1395 = mem_3[tmp1220];
    assign tmp2554 = {tmp2553[0], tmp2553[1], tmp2553[2], tmp2553[3], tmp2553[4], tmp2553[5], tmp2553[6], tmp2553[7]};
    assign tmp2407 = tmp2566;
        assign tmp2350 = mem_1[tmp2318];
    assign b4_w7 = tmp42;
    assign tmp2575 = {const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0, const2574_0};
    assign tmp1425 = tmp1421 ^ tmp1424;
        assign tmp1472 = mem_1[tmp1440];
    assign tmp1409 = tmp1407 ^ tmp1408;
    assign tmp1657 = {tmp1656, tmp1508};
    assign tmp576 = tmp592;
    assign tmp2833 = {tmp2832, tmp2681};
    assign tmp2499 = {const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0, const2498_0};
    assign rc2_w15 = const100_0;
    assign c2_w39 = tmp244;
    assign tmp2417 = tmp2413 ^ tmp2416;
    assign tmp324 = {temp_1[16], temp_1[17], temp_1[18], temp_1[19], temp_1[20], temp_1[21], temp_1[22], temp_1[23]};
        assign tmp834 = mem_4[tmp633];
    assign tmp2726 = tmp2722 ^ tmp2725;
        assign tmp713 = mem_3[tmp626];
    assign tmp2929 = tmp2945;
    assign tmp1368 = {tmp1367, tmp1216};
    assign tmp2047 = tmp2063;
    assign tmp802 = {tmp801, tmp635};
    assign tmp2621 = {temp_32[0], temp_32[1], temp_32[2], temp_32[3], temp_32[4], temp_32[5], temp_32[6], temp_32[7]};
    assign tmp927 = {temp_10[16], temp_10[17], temp_10[18], temp_10[19], temp_10[20], temp_10[21], temp_10[22], temp_10[23]};
        assign tmp786 = mem_4[tmp629];
    assign tmp2088 = {temp_26[104], temp_26[105], temp_26[106], temp_26[107], temp_26[108], temp_26[109], temp_26[110], temp_26[111]};
    assign tmp581 = tmp597;
    assign shifted_w39 = tmp238;
    assign tmp2834 = tmp2830 ^ tmp2833;
        assign tmp1665 = mem_4[tmp1508];
    assign tmp2032 = {temp_24[24], temp_24[25], temp_24[26], temp_24[27], temp_24[28], temp_24[29], temp_24[30], temp_24[31]};
    assign tmp644 = tmp748;
        assign tmp2753 = mem_4[tmp2677];
    assign tmp2444 = {tmp2443, tmp2380};
    assign tmp603 = {tmp571, tmp572, tmp573, tmp574, tmp575, tmp576, tmp577, tmp578, tmp579, tmp580, tmp581, tmp582, tmp583, tmp584, tmp585, tmp586};
        assign tmp1067 = mem_4[tmp925];
    assign tmp2323 = {temp_28[40], temp_28[41], temp_28[42], temp_28[43], temp_28[44], temp_28[45], temp_28[46], temp_28[47]};
        assign tmp1580 = mem_3[tmp1504];
    assign tmp2017 = {tmp1809, tmp1810, tmp1811, tmp1812, tmp1813, tmp1814, tmp1815, tmp1816, tmp1817, tmp1818, tmp1819, tmp1820, tmp1821, tmp1822, tmp1823, tmp1824};
    assign tmp1144 = {temp_12[96], temp_12[97], temp_12[98], temp_12[99], temp_12[100], temp_12[101], temp_12[102], temp_12[103]};
    assign shifted_w23 = tmp138;
        assign tmp145 = mem_1[b3_w23];
        assign tmp1360 = mem_4[tmp1218];
    assign tmp1783 = {temp_21[64], temp_21[65], temp_21[66], temp_21[67], temp_21[68], temp_21[69], temp_21[70], temp_21[71]};
        assign tmp1384 = mem_4[tmp1220];
    assign tmp1681 = {tmp1680, tmp1514};
    assign tmp796 = {tmp795[0], tmp795[1], tmp795[2], tmp795[3], tmp795[4], tmp795[5], tmp795[6], tmp795[7]};
    assign substituted_w31 = tmp197;
    assign tmp1866 = {tmp1865, tmp1794};
    assign tmp270 = {new_state[56], new_state[57], new_state[58], new_state[59], new_state[60], new_state[61], new_state[62], new_state[63]};
    assign tmp1459 = tmp1475;
    assign tmp1071 = {tmp1070, tmp922};
    assign tmp1041 = {tmp1040[0], tmp1040[1], tmp1040[2], tmp1040[3], tmp1040[4], tmp1040[5], tmp1040[6], tmp1040[7]};
    assign tmp2693 = tmp2775;
    assign tmp1555 = {tmp1554[0], tmp1554[1], tmp1554[2], tmp1554[3], tmp1554[4], tmp1554[5], tmp1554[6], tmp1554[7]};
    assign tmp1602 = tmp1598 ^ tmp1601;
    assign tmp2101 = {temp_26[0], temp_26[1], temp_26[2], temp_26[3], temp_26[4], temp_26[5], temp_26[6], temp_26[7]};
    assign tmp2866 = tmp2862 ^ tmp2865;
    assign tmp2718 = tmp2716 ^ tmp2717;
    assign tmp496 = {const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0, const495_0};
    assign tmp458 = tmp456 ^ tmp457;
        assign tmp1407 = mem_3[tmp1221];
    assign tmp978 = {const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0, const977_0};
    assign tmp1428 = {tmp1427, tmp1221};
        assign tmp2643 = mem_1[tmp2611];
    assign tmp2919 = tmp2935;
    assign tmp1717 = {tmp1716, tmp1513};
    assign tmp562 = {temp_4[64], temp_4[65], temp_4[66], temp_4[67], temp_4[68], temp_4[69], temp_4[70], temp_4[71]};
    assign new_2 = tmp554;
    assign tmp242 = {shifted_w39[0], shifted_w39[1], shifted_w39[2], shifted_w39[3], shifted_w39[4], shifted_w39[5], shifted_w39[6], shifted_w39[7]};
    assign tmp141 = {shifted_w23[8], shifted_w23[9], shifted_w23[10], shifted_w23[11], shifted_w23[12], shifted_w23[13], shifted_w23[14], shifted_w23[15]};
    assign tmp921 = {temp_10[64], temp_10[65], temp_10[66], temp_10[67], temp_10[68], temp_10[69], temp_10[70], temp_10[71]};
        assign tmp2356 = mem_1[tmp2324];
    assign tmp1022 = {const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0, const1021_0};
    assign a4_w35 = tmp212;
    assign tmp2713 = {tmp2712, tmp2675};
        assign tmp2825 = mem_4[tmp2683];
    assign tmp897 = {temp_9[120], temp_9[121], temp_9[122], temp_9[123], temp_9[124], temp_9[125], temp_9[126], temp_9[127]};
    assign temp_26 = tmp2085;
    assign tmp2668 = {temp_33[16], temp_33[17], temp_33[18], temp_33[19], temp_33[20], temp_33[21], temp_33[22], temp_33[23]};
    assign tmp2667 = {temp_33[24], temp_33[25], temp_33[26], temp_33[27], temp_33[28], temp_33[29], temp_33[30], temp_33[31]};
    assign tmp321 = {temp_1[40], temp_1[41], temp_1[42], temp_1[43], temp_1[44], temp_1[45], temp_1[46], temp_1[47]};
    assign a3_w19 = tmp111;
    assign c1_w19 = tmp118;
    assign tmp682 = {tmp681, tmp621};
        assign tmp1771 = mem_1[tmp1739];
    assign tmp1397 = tmp1395 ^ tmp1396;
        assign tmp1078 = mem_3[tmp925];
    assign tmp1615 = {tmp1614[0], tmp1614[1], tmp1614[2], tmp1614[3], tmp1614[4], tmp1614[5], tmp1614[6], tmp1614[7]};
    assign tmp2894 = tmp2890 ^ tmp2893;
    assign tmp1423 = {const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0, const1422_0};
    assign tmp2802 = tmp2800 ^ tmp2801;
        assign tmp1030 = mem_3[tmp921];
    assign tmp2075 = {temp_25[72], temp_25[73], temp_25[74], temp_25[75], temp_25[76], temp_25[77], temp_25[78], temp_25[79]};
        assign tmp1994 = mem_4[tmp1808];
        assign tmp169 = mem_1[b2_w27];
    assign tmp2441 = tmp2437 ^ tmp2440;
        assign tmp1886 = mem_4[tmp1799];
        assign tmp2215 = mem_4[tmp2095];
    assign tmp2416 = {tmp2415, tmp2381};
    assign tmp1134 = {const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0, const1133_0};
    assign tmp1245 = tmp1241 ^ tmp1244;
        assign tmp590 = mem_1[tmp558];
    assign tmp2916 = tmp2932;
    assign tmp2335 = tmp2351;
        assign tmp2411 = mem_3[tmp2379];
        assign tmp1569 = mem_4[tmp1500];
    assign tmp2908 = {temp_36[48], temp_36[49], temp_36[50], temp_36[51], temp_36[52], temp_36[53], temp_36[54], temp_36[55]};
    assign tmp1322 = {tmp1321[0], tmp1321[1], tmp1321[2], tmp1321[3], tmp1321[4], tmp1321[5], tmp1321[6], tmp1321[7]};
    assign tmp2537 = tmp2533 ^ tmp2536;
    assign tmp253 = {rc1_w39, rc2_w39, rc3_w39, rc4_w39};
    assign tmp926 = {temp_10[24], temp_10[25], temp_10[26], temp_10[27], temp_10[28], temp_10[29], temp_10[30], temp_10[31]};
    assign tmp857 = {temp_8[48], temp_8[49], temp_8[50], temp_8[51], temp_8[52], temp_8[53], temp_8[54], temp_8[55]};
    assign tmp2781 = {tmp2780, tmp2676};
        assign tmp1371 = mem_3[tmp1218];
    assign tmp2162 = {const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0, const2161_0};
    assign tmp2610 = {temp_32[88], temp_32[89], temp_32[90], temp_32[91], temp_32[92], temp_32[93], temp_32[94], temp_32[95]};
        assign tmp480 = mem_3[tmp338];
    assign tmp2511 = {const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0, const2510_0};
        assign tmp2642 = mem_1[tmp2610];
    assign tmp582 = tmp598;
    assign tmp1147 = {temp_12[72], temp_12[73], temp_12[74], temp_12[75], temp_12[76], temp_12[77], temp_12[78], temp_12[79]};
    assign tmp2625 = tmp2641;
    assign tmp1638 = tmp1634 ^ tmp1637;
    assign tmp1990 = {tmp1989, tmp1805};
    assign tmp2778 = tmp2776 ^ tmp2777;
        assign tmp309 = mem_1[tmp277];
    assign tmp908 = {temp_9[32], temp_9[33], temp_9[34], temp_9[35], temp_9[36], temp_9[37], temp_9[38], temp_9[39]};
        assign tmp294 = mem_1[tmp262];
    assign tmp2614 = {temp_32[56], temp_32[57], temp_32[58], temp_32[59], temp_32[60], temp_32[61], temp_32[62], temp_32[63]};
    assign tmp1044 = tmp1042 ^ tmp1043;
    assign tmp952 = tmp948 ^ tmp951;
    assign tmp2292 = tmp2288 ^ tmp2291;
    assign tmp650 = tmp820;
    assign tmp734 = {tmp733, tmp626};
    assign tmp984 = tmp982 ^ tmp983;
    assign tmp1393 = tmp1389 ^ tmp1392;
    assign tmp2489 = tmp2485 ^ tmp2488;
    assign tmp1807 = {temp_22[8], temp_22[9], temp_22[10], temp_22[11], temp_22[12], temp_22[13], temp_22[14], temp_22[15]};
    assign tmp1504 = {temp_18[88], temp_18[89], temp_18[90], temp_18[91], temp_18[92], temp_18[93], temp_18[94], temp_18[95]};
    assign tmp2515 = {const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0, const2514_0};
    assign tmp2267 = {tmp2266, tmp2100};
    assign tmp1026 = {const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0, const1025_0};
    assign tmp2862 = tmp2860 ^ tmp2861;
    assign tmp353 = tmp479;
    assign tmp1870 = {tmp1869, tmp1795};
    assign tmp1997 = {const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0, const1996_0};
    assign a2_w15 = tmp85;
        assign tmp2496 = mem_4[tmp2383];
    assign tmp1135 = {tmp1134, tmp928};
    assign tmp2859 = {tmp2858[0], tmp2858[1], tmp2858[2], tmp2858[3], tmp2858[4], tmp2858[5], tmp2858[6], tmp2858[7]};
    assign temp_7 = tmp845;
    assign tmp585 = tmp601;
    assign tmp975 = {tmp974, tmp914};
    assign tmp1596 = {const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0, const1595_0};
    assign tmp1232 = tmp1358;
    assign substituted_w35 = tmp222;
    assign tmp1358 = {tmp1357[0], tmp1357[1], tmp1357[2], tmp1357[3], tmp1357[4], tmp1357[5], tmp1357[6], tmp1357[7]};
    assign c4_w35 = tmp221;
    assign tmp1280 = {tmp1279, tmp1208};
    assign tmp625 = {temp_6[88], temp_6[89], temp_6[90], temp_6[91], temp_6[92], temp_6[93], temp_6[94], temp_6[95]};
        assign tmp1713 = mem_4[tmp1512];
    assign tmp769 = {const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0, const768_0};
    assign tmp2923 = tmp2939;
    assign tmp967 = {tmp966, tmp914};
        assign tmp601 = mem_1[tmp569];
        assign tmp195 = mem_1[b3_w31];
    assign tmp1464 = tmp1480;
    assign rc2_w39 = const250_0;
    assign c3_w35 = tmp220;
    assign tmp1877 = {const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0, const1876_0};
    assign tmp1847 = tmp1843 ^ tmp1846;
    assign tmp1646 = tmp1642 ^ tmp1645;
    assign tmp1558 = tmp1556 ^ tmp1557;
        assign tmp2142 = mem_3[tmp2088];
    assign concat_w19 = tmp128;
    assign tmp1400 = {tmp1399, tmp1222};
    assign tmp758 = {tmp757, tmp632};
    assign tmp1435 = {temp_16[112], temp_16[113], temp_16[114], temp_16[115], temp_16[116], temp_16[117], temp_16[118], temp_16[119]};
    assign tmp1987 = tmp1983 ^ tmp1986;
    assign tmp2602 = {tmp2601[0], tmp2601[1], tmp2601[2], tmp2601[3], tmp2601[4], tmp2601[5], tmp2601[6], tmp2601[7]};
    assign tmp2549 = tmp2545 ^ tmp2548;
    assign tmp382 = tmp378 ^ tmp381;
    assign tmp1649 = {tmp1648, tmp1508};
    assign tmp1098 = {const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0, const1097_0};
    assign tmp1514 = {temp_18[8], temp_18[9], temp_18[10], temp_18[11], temp_18[12], temp_18[13], temp_18[14], temp_18[15]};
    assign shifted_w31 = tmp188;
    assign tmp28 = {rc1_w3, rc2_w3, rc3_w3, rc4_w3};
        assign tmp120 = mem_1[b3_w19];
    assign tmp359 = tmp551;
    assign tmp1027 = {tmp1026, tmp919};
    assign tmp1780 = {temp_21[88], temp_21[89], temp_21[90], temp_21[91], temp_21[92], temp_21[93], temp_21[94], temp_21[95]};
    assign tmp422 = tmp420 ^ tmp421;
        assign tmp2946 = mem_1[tmp2914];
    assign tmp33 = w6 ^ w3;
    assign tmp1734 = {temp_20[64], temp_20[65], temp_20[66], temp_20[67], temp_20[68], temp_20[69], temp_20[70], temp_20[71]};
    assign a4_w11 = tmp62;
    assign tmp2433 = tmp2429 ^ tmp2432;
    assign concat_w27 = tmp178;
    assign tmp830 = {tmp829, tmp634};
    assign tmp35 = {w7[16], w7[17], w7[18], w7[19], w7[20], w7[21], w7[22], w7[23]};
    assign tmp2041 = tmp2057;
        assign tmp2935 = mem_1[tmp2903];
    assign a4_w7 = tmp37;
    assign tmp730 = {tmp729, tmp625};
    assign tmp1227 = tmp1298;
    assign tmp2672 = {temp_34[120], temp_34[121], temp_34[122], temp_34[123], temp_34[124], temp_34[125], temp_34[126], temp_34[127]};
    assign tmp1507 = {temp_18[64], temp_18[65], temp_18[66], temp_18[67], temp_18[68], temp_18[69], temp_18[70], temp_18[71]};
    assign tmp1110 = {const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0, const1109_0};
    assign tmp2868 = {const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0, const2867_0};
    assign a2_w23 = tmp135;
    assign tmp782 = {tmp781, tmp630};
        assign tmp2788 = mem_3[tmp2679];
    assign c1_w23 = tmp143;
    assign tmp502 = tmp498 ^ tmp501;
    assign tmp526 = tmp522 ^ tmp525;
    assign tmp1823 = tmp2004;
        assign tmp1481 = mem_1[tmp1449];
    assign tmp2627 = tmp2643;
    assign tmp2584 = {tmp2583, tmp2391};
    assign tmp2733 = {tmp2732, tmp2672};
    assign tmp1198 = {temp_13[56], temp_13[57], temp_13[58], temp_13[59], temp_13[60], temp_13[61], temp_13[62], temp_13[63]};
    assign b4_w27 = tmp167;
        assign tmp690 = mem_4[tmp621];
    assign tmp1197 = {temp_13[64], temp_13[65], temp_13[66], temp_13[67], temp_13[68], temp_13[69], temp_13[70], temp_13[71]};
    assign concat_w7 = tmp53;
    assign tmp900 = {temp_9[96], temp_9[97], temp_9[98], temp_9[99], temp_9[100], temp_9[101], temp_9[102], temp_9[103]};
        assign tmp2740 = mem_3[tmp2675];
    assign tmp2512 = {tmp2511, tmp2389};
        assign tmp1910 = mem_4[tmp1797];
    assign tmp277 = {new_state[0], new_state[1], new_state[2], new_state[3], new_state[4], new_state[5], new_state[6], new_state[7]};
    assign tmp328 = {temp_2[120], temp_2[121], temp_2[122], temp_2[123], temp_2[124], temp_2[125], temp_2[126], temp_2[127]};
    assign tmp2039 = tmp2055;
    assign tmp1606 = tmp1604 ^ tmp1605;
        assign tmp892 = mem_1[tmp860];
        assign tmp1006 = mem_3[tmp919];
    assign tmp1172 = tmp1188;
    assign rc4_w31 = const202_0;
    assign tmp1621 = {tmp1620, tmp1505};
    assign tmp979 = {tmp978, tmp915};
    assign tmp2521 = tmp2519 ^ tmp2520;
        assign tmp2520 = mem_4[tmp2389];
        assign tmp2519 = mem_3[tmp2388];
    assign w1 = tmp6;
        assign tmp2789 = mem_4[tmp2676];
    assign tmp845 = {tmp637, tmp638, tmp639, tmp640, tmp641, tmp642, tmp643, tmp644, tmp645, tmp646, tmp647, tmp648, tmp649, tmp650, tmp651, tmp652};
    assign tmp2319 = {temp_28[72], temp_28[73], temp_28[74], temp_28[75], temp_28[76], temp_28[77], temp_28[78], temp_28[79]};
    assign tmp2314 = {temp_28[112], temp_28[113], temp_28[114], temp_28[115], temp_28[116], temp_28[117], temp_28[118], temp_28[119]};
        assign tmp1476 = mem_1[tmp1444];
        assign tmp2460 = mem_4[tmp2384];
    assign tmp1403 = {const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0, const1402_0};
    assign tmp181 = tmp180 ^ tmp156;
    assign tmp1141 = {temp_12[120], temp_12[121], temp_12[122], temp_12[123], temp_12[124], temp_12[125], temp_12[126], temp_12[127]};
        assign tmp302 = mem_1[tmp270];
    assign tmp1790 = {temp_21[8], temp_21[9], temp_21[10], temp_21[11], temp_21[12], temp_21[13], temp_21[14], temp_21[15]};
    assign tmp42 = {shifted_w7[0], shifted_w7[1], shifted_w7[2], shifted_w7[3], shifted_w7[4], shifted_w7[5], shifted_w7[6], shifted_w7[7]};
    assign tmp278 = tmp294;
    assign tmp2589 = tmp2585 ^ tmp2588;
    assign tmp2182 = {const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0, const2181_0};
    assign tmp2216 = tmp2214 ^ tmp2215;
    assign tmp2288 = tmp2286 ^ tmp2287;
    assign tmp1716 = {const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0, const1715_0};
        assign tmp1766 = mem_1[tmp1734];
    assign tmp414 = tmp410 ^ tmp413;
    assign tmp1375 = {const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0, const1374_0};
    assign tmp2809 = {tmp2808, tmp2683};
    assign tmp135 = {tmp133[16], tmp133[17], tmp133[18], tmp133[19], tmp133[20], tmp133[21], tmp133[22], tmp133[23]};
    assign tmp247 = {c1_w39, c2_w39, c3_w39, c4_w39};
    assign tmp1216 = {temp_14[48], temp_14[49], temp_14[50], temp_14[51], temp_14[52], temp_14[53], temp_14[54], temp_14[55]};
    assign w3 = tmp8;
    assign tmp233 = tmp232 ^ tmp208;
    assign tmp2787 = {tmp2786[0], tmp2786[1], tmp2786[2], tmp2786[3], tmp2786[4], tmp2786[5], tmp2786[6], tmp2786[7]};
    assign tmp89 = {shifted_w15[24], shifted_w15[25], shifted_w15[26], shifted_w15[27], shifted_w15[28], shifted_w15[29], shifted_w15[30], shifted_w15[31]};
        assign tmp492 = mem_3[tmp339];
    assign tmp1279 = {const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0, const1278_0};
    assign tmp2300 = tmp2298 ^ tmp2299;
        assign tmp1102 = mem_3[tmp927];
    assign tmp1782 = {temp_21[72], temp_21[73], temp_21[74], temp_21[75], temp_21[76], temp_21[77], temp_21[78], temp_21[79]};
    assign tmp938 = tmp1053;
        assign tmp2483 = mem_3[tmp2385];
    assign tmp2174 = {const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0, const2173_0};
    assign tmp1052 = tmp1048 ^ tmp1051;
        assign tmp168 = mem_1[b1_w27];
    assign tmp2107 = tmp2189;
    assign tmp2027 = {temp_24[64], temp_24[65], temp_24[66], temp_24[67], temp_24[68], temp_24[69], temp_24[70], temp_24[71]};
    assign tmp2050 = tmp2066;
    assign tmp2950 = {temp_37[104], temp_37[105], temp_37[106], temp_37[107], temp_37[108], temp_37[109], temp_37[110], temp_37[111]};
    assign tmp1540 = {const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0, const1539_0};
    assign tmp38 = {a2_w7, a3_w7, a4_w7, a1_w7};
        assign tmp2061 = mem_1[tmp2029];
    assign tmp1377 = tmp1373 ^ tmp1376;
    assign c1_w7 = tmp43;
        assign tmp2154 = mem_3[tmp2089];
        assign tmp95 = mem_1[b3_w15];
    assign tmp2463 = {const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0, const2462_0};
    assign tmp1367 = {const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0, const1366_0};
    assign tmp757 = {const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0, const756_0};
    assign tmp1332 = {tmp1331, tmp1213};
    assign tmp2684 = {temp_34[24], temp_34[25], temp_34[26], temp_34[27], temp_34[28], temp_34[29], temp_34[30], temp_34[31]};
    assign tmp2051 = tmp2067;
    assign tmp1867 = tmp1863 ^ tmp1866;
    assign tmp1125 = {tmp1124[0], tmp1124[1], tmp1124[2], tmp1124[3], tmp1124[4], tmp1124[5], tmp1124[6], tmp1124[7]};
    assign tmp2406 = tmp2554;
    assign tmp2664 = {temp_33[48], temp_33[49], temp_33[50], temp_33[51], temp_33[52], temp_33[53], temp_33[54], temp_33[55]};
    assign tmp430 = tmp426 ^ tmp429;
    assign tmp449 = {tmp448, tmp333};
    assign tmp1234 = tmp1382;
    assign tmp1017 = {tmp1016[0], tmp1016[1], tmp1016[2], tmp1016[3], tmp1016[4], tmp1016[5], tmp1016[6], tmp1016[7]};
    assign tmp1577 = {tmp1576, tmp1502};
    assign tmp64 = {shifted_w11[24], shifted_w11[25], shifted_w11[26], shifted_w11[27], shifted_w11[28], shifted_w11[29], shifted_w11[30], shifted_w11[31]};
    assign tmp1903 = tmp1899 ^ tmp1902;
    assign tmp390 = tmp386 ^ tmp389;
    assign tmp216 = {shifted_w35[8], shifted_w35[9], shifted_w35[10], shifted_w35[11], shifted_w35[12], shifted_w35[13], shifted_w35[14], shifted_w35[15]};
        assign tmp678 = mem_4[tmp624];
        assign tmp2435 = mem_3[tmp2381];
    assign tmp1148 = {temp_12[64], temp_12[65], temp_12[66], temp_12[67], temp_12[68], temp_12[69], temp_12[70], temp_12[71]};
    assign tmp47 = {c1_w7, c2_w7, c3_w7, c4_w7};
    assign tmp2692 = tmp2763;
    assign tmp966 = {const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0, const965_0};
    assign tmp548 = {const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0, const547_0};
        assign tmp303 = mem_1[tmp271];
    assign tmp808 = {tmp807[0], tmp807[1], tmp807[2], tmp807[3], tmp807[4], tmp807[5], tmp807[6], tmp807[7]};
    assign tmp90 = {shifted_w15[16], shifted_w15[17], shifted_w15[18], shifted_w15[19], shifted_w15[20], shifted_w15[21], shifted_w15[22], shifted_w15[23]};
        assign tmp891 = mem_1[tmp859];
    assign tmp1482 = {tmp1450, tmp1451, tmp1452, tmp1453, tmp1454, tmp1455, tmp1456, tmp1457, tmp1458, tmp1459, tmp1460, tmp1461, tmp1462, tmp1463, tmp1464, tmp1465};
    assign tmp2636 = tmp2652;
    assign tmp1165 = tmp1181;
        assign tmp1466 = mem_1[tmp1434];
    assign tmp806 = {tmp805, tmp636};
        assign tmp1335 = mem_3[tmp1215];
    assign tmp1699 = {tmp1698[0], tmp1698[1], tmp1698[2], tmp1698[3], tmp1698[4], tmp1698[5], tmp1698[6], tmp1698[7]};
        assign tmp959 = mem_4[tmp916];
    assign tmp2153 = {tmp2152[0], tmp2152[1], tmp2152[2], tmp2152[3], tmp2152[4], tmp2152[5], tmp2152[6], tmp2152[7]};
    assign tmp1153 = {temp_12[24], temp_12[25], temp_12[26], temp_12[27], temp_12[28], temp_12[29], temp_12[30], temp_12[31]};
    assign tmp211 = {tmp208[8], tmp208[9], tmp208[10], tmp208[11], tmp208[12], tmp208[13], tmp208[14], tmp208[15]};
    assign rc1_w7 = tmp49;
        assign tmp994 = mem_3[tmp918];
    assign tmp1190 = {temp_13[120], temp_13[121], temp_13[122], temp_13[123], temp_13[124], temp_13[125], temp_13[126], temp_13[127]};
    assign a2_w19 = tmp110;
    assign tmp2844 = {const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0, const2843_0};
    assign tmp344 = tmp371;
    assign new_3 = tmp847;
    assign tmp443 = {tmp442[0], tmp442[1], tmp442[2], tmp442[3], tmp442[4], tmp442[5], tmp442[6], tmp442[7]};
        assign tmp882 = mem_1[tmp850];
    assign aes_ciphertext = temp_39;
        assign tmp174 = mem_2[const173_7];
    assign tmp765 = {const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0, const764_0};
    assign tmp663 = tmp659 ^ tmp662;
    assign tmp1741 = {temp_20[8], temp_20[9], temp_20[10], temp_20[11], temp_20[12], temp_20[13], temp_20[14], temp_20[15]};
        assign tmp1183 = mem_1[tmp1151];
    assign tmp1935 = tmp1933 ^ tmp1934;
    assign tmp2703 = tmp2895;
    assign tmp407 = {tmp406[0], tmp406[1], tmp406[2], tmp406[3], tmp406[4], tmp406[5], tmp406[6], tmp406[7]};
    assign tmp913 = {tmp897, tmp902, tmp907, tmp912, tmp901, tmp906, tmp911, tmp900, tmp905, tmp910, tmp899, tmp904, tmp909, tmp898, tmp903, tmp908};
    assign tmp2388 = {temp_30[48], temp_30[49], temp_30[50], temp_30[51], temp_30[52], temp_30[53], temp_30[54], temp_30[55]};
    assign tmp699 = tmp695 ^ tmp698;
    assign tmp1798 = {temp_22[80], temp_22[81], temp_22[82], temp_22[83], temp_22[84], temp_22[85], temp_22[86], temp_22[87]};
    assign tmp317 = {temp_1[72], temp_1[73], temp_1[74], temp_1[75], temp_1[76], temp_1[77], temp_1[78], temp_1[79]};
        assign tmp1312 = mem_4[tmp1214];
    assign tmp742 = {tmp741, tmp626};
        assign tmp2355 = mem_1[tmp2323];
        assign tmp2238 = mem_3[tmp2096];
    assign shifted_w19 = tmp113;
        assign tmp1477 = mem_1[tmp1445];
    assign tmp1854 = {tmp1853, tmp1793};
    assign tmp157 = tmp156 ^ tmp132;
    assign rc3_w7 = const51_0;
        assign tmp2716 = mem_3[tmp2673];
    assign tmp2270 = {const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0, const2269_0};
    assign tmp2656 = {temp_33[112], temp_33[113], temp_33[114], temp_33[115], temp_33[116], temp_33[117], temp_33[118], temp_33[119]};
    assign temp_31 = tmp2603;
    assign tmp257 = tmp256 ^ tmp232;
    assign tmp2749 = {tmp2748, tmp2674};
        assign tmp2348 = mem_1[tmp2316];
    assign a2_w31 = tmp185;
    assign rc3_w11 = const76_0;
    assign tmp1711 = {tmp1710[0], tmp1710[1], tmp1710[2], tmp1710[3], tmp1710[4], tmp1710[5], tmp1710[6], tmp1710[7]};
    assign tmp1746 = tmp1762;
    assign tmp2780 = {const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0, const2779_0};
        assign tmp1467 = mem_1[tmp1435];
    assign input_wire_3 = temp_7;
    assign tmp2186 = {const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0, const2185_0};
    assign tmp2654 = {tmp2622, tmp2623, tmp2624, tmp2625, tmp2626, tmp2627, tmp2628, tmp2629, tmp2630, tmp2631, tmp2632, tmp2633, tmp2634, tmp2635, tmp2636, tmp2637};
    assign tmp1461 = tmp1477;
    assign tmp1131 = {tmp1130, tmp927};
    assign tmp1818 = tmp1944;
        assign tmp2934 = mem_1[tmp2902];
    assign tmp1099 = {tmp1098, tmp929};
    assign tmp2766 = tmp2764 ^ tmp2765;
    assign tmp729 = {const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0, const728_0};
    assign tmp826 = {tmp825, tmp633};
    assign tmp1490 = {temp_17[64], temp_17[65], temp_17[66], temp_17[67], temp_17[68], temp_17[69], temp_17[70], temp_17[71]};
    assign b1_w27 = tmp164;
    assign tmp203 = {rc1_w31, rc2_w31, rc3_w31, rc4_w31};
        assign tmp592 = mem_1[tmp560];
    assign tmp2925 = tmp2941;
    assign tmp1673 = {tmp1672, tmp1510};
    assign tmp406 = tmp402 ^ tmp405;
    assign tmp2261 = {tmp2260[0], tmp2260[1], tmp2260[2], tmp2260[3], tmp2260[4], tmp2260[5], tmp2260[6], tmp2260[7]};
    assign tmp1610 = tmp1606 ^ tmp1609;
    assign tmp2898 = temp_35 ^ tmp2897;
    assign tmp1656 = {const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0, const1655_0};
    assign tmp1857 = {const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0, const1856_0};
    assign tmp956 = tmp952 ^ tmp955;
        assign tmp2938 = mem_1[tmp2906];
    assign tmp2961 = {temp_37[16], temp_37[17], temp_37[18], temp_37[19], temp_37[20], temp_37[21], temp_37[22], temp_37[23]};
    assign a1_w19 = tmp109;
        assign tmp296 = mem_1[tmp264];
    assign tmp681 = {const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0, const680_0};
        assign tmp1629 = mem_4[tmp1509];
        assign tmp1861 = mem_3[tmp1796];
    assign tmp2810 = tmp2806 ^ tmp2809;
    assign tmp1196 = {temp_13[72], temp_13[73], temp_13[74], temp_13[75], temp_13[76], temp_13[77], temp_13[78], temp_13[79]};
    assign tmp155 = tmp130 ^ xor_w23;
    assign tmp1496 = {temp_17[16], temp_17[17], temp_17[18], temp_17[19], temp_17[20], temp_17[21], temp_17[22], temp_17[23]};
    assign temp_12 = new_4;
        assign tmp889 = mem_1[tmp857];
    assign tmp2604 = {expanded_key[256], expanded_key[257], expanded_key[258], expanded_key[259], expanded_key[260], expanded_key[261], expanded_key[262], expanded_key[263], expanded_key[264], expanded_key[265], expanded_key[266], expanded_key[267], expanded_key[268], expanded_key[269], expanded_key[270], expanded_key[271], expanded_key[272], expanded_key[273], expanded_key[274], expanded_key[275], expanded_key[276], expanded_key[277], expanded_key[278], expanded_key[279], expanded_key[280], expanded_key[281], expanded_key[282], expanded_key[283], expanded_key[284], expanded_key[285], expanded_key[286], expanded_key[287], expanded_key[288], expanded_key[289], expanded_key[290], expanded_key[291], expanded_key[292], expanded_key[293], expanded_key[294], expanded_key[295], expanded_key[296], expanded_key[297], expanded_key[298], expanded_key[299], expanded_key[300], expanded_key[301], expanded_key[302], expanded_key[303], expanded_key[304], expanded_key[305], expanded_key[306], expanded_key[307], expanded_key[308], expanded_key[309], expanded_key[310], expanded_key[311], expanded_key[312], expanded_key[313], expanded_key[314], expanded_key[315], expanded_key[316], expanded_key[317], expanded_key[318], expanded_key[319], expanded_key[320], expanded_key[321], expanded_key[322], expanded_key[323], expanded_key[324], expanded_key[325], expanded_key[326], expanded_key[327], expanded_key[328], expanded_key[329], expanded_key[330], expanded_key[331], expanded_key[332], expanded_key[333], expanded_key[334], expanded_key[335], expanded_key[336], expanded_key[337], expanded_key[338], expanded_key[339], expanded_key[340], expanded_key[341], expanded_key[342], expanded_key[343], expanded_key[344], expanded_key[345], expanded_key[346], expanded_key[347], expanded_key[348], expanded_key[349], expanded_key[350], expanded_key[351], expanded_key[352], expanded_key[353], expanded_key[354], expanded_key[355], expanded_key[356], expanded_key[357], expanded_key[358], expanded_key[359], expanded_key[360], expanded_key[361], expanded_key[362], expanded_key[363], expanded_key[364], expanded_key[365], expanded_key[366], expanded_key[367], expanded_key[368], expanded_key[369], expanded_key[370], expanded_key[371], expanded_key[372], expanded_key[373], expanded_key[374], expanded_key[375], expanded_key[376], expanded_key[377], expanded_key[378], expanded_key[379], expanded_key[380], expanded_key[381], expanded_key[382], expanded_key[383]};
        assign tmp2531 = mem_3[tmp2389];
    assign tmp1303 = {const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0, const1302_0};
    assign tmp2105 = tmp2165;
    assign tmp1363 = {const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0, const1362_0};
    assign tmp1456 = tmp1472;
    assign tmp2310 = {tmp2102, tmp2103, tmp2104, tmp2105, tmp2106, tmp2107, tmp2108, tmp2109, tmp2110, tmp2111, tmp2112, tmp2113, tmp2114, tmp2115, tmp2116, tmp2117};
    assign tmp2737 = {tmp2736, tmp2673};
    assign tmp627 = {temp_6[72], temp_6[73], temp_6[74], temp_6[75], temp_6[76], temp_6[77], temp_6[78], temp_6[79]};
    assign tmp827 = tmp823 ^ tmp826;
    assign tmp741 = {const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0, const740_0};
    assign tmp2663 = {temp_33[56], temp_33[57], temp_33[58], temp_33[59], temp_33[60], temp_33[61], temp_33[62], temp_33[63]};
    assign rc2_w7 = const50_0;
    assign tmp2211 = {tmp2210, tmp2092};
    assign tmp2093 = {temp_26[64], temp_26[65], temp_26[66], temp_26[67], temp_26[68], temp_26[69], temp_26[70], temp_26[71]};
    assign tmp2870 = tmp2866 ^ tmp2869;
    assign tmp153 = {rc1_w23, rc2_w23, rc3_w23, rc4_w23};
    assign tmp1816 = tmp1920;
    assign tmp85 = {tmp83[16], tmp83[17], tmp83[18], tmp83[19], tmp83[20], tmp83[21], tmp83[22], tmp83[23]};
    assign tmp138 = {a2_w23, a3_w23, a4_w23, a1_w23};
    assign tmp342 = {temp_2[8], temp_2[9], temp_2[10], temp_2[11], temp_2[12], temp_2[13], temp_2[14], temp_2[15]};
    assign tmp2701 = tmp2871;
        assign tmp372 = mem_3[tmp329];
    assign tmp186 = {tmp183[8], tmp183[9], tmp183[10], tmp183[11], tmp183[12], tmp183[13], tmp183[14], tmp183[15]};
    assign tmp1710 = tmp1706 ^ tmp1709;
    assign tmp1231 = tmp1346;
        assign tmp982 = mem_3[tmp917];
    assign tmp1271 = {const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0, const1270_0};
    assign tmp370 = tmp366 ^ tmp369;
    assign tmp1588 = {const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0, const1587_0};
    assign a3_w39 = tmp236;
    assign tmp398 = tmp396 ^ tmp397;
    assign tmp2905 = {temp_36[72], temp_36[73], temp_36[74], temp_36[75], temp_36[76], temp_36[77], temp_36[78], temp_36[79]};
        assign tmp1103 = mem_4[tmp928];
        assign tmp74 = mem_2[const73_3];
        assign tmp1767 = mem_1[tmp1735];
    assign tmp1967 = tmp1963 ^ tmp1966;
    assign tmp425 = {tmp424, tmp335};
    assign tmp1723 = {tmp1722[0], tmp1722[1], tmp1722[2], tmp1722[3], tmp1722[4], tmp1722[5], tmp1722[6], tmp1722[7]};
    assign tmp1651 = {tmp1650[0], tmp1650[1], tmp1650[2], tmp1650[3], tmp1650[4], tmp1650[5], tmp1650[6], tmp1650[7]};
    assign temp_10 = tmp913;
    assign tmp2246 = {const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0, const2245_0};
    assign tmp831 = tmp827 ^ tmp830;
    assign tmp1930 = {tmp1929, tmp1804};
    assign tmp2551 = {const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0, const2550_0};
    assign tmp2881 = {tmp2880, tmp2685};
    assign tmp287 = tmp303;
        assign tmp384 = mem_3[tmp330];
    assign tmp1726 = temp_19 ^ tmp1725;
    assign tmp346 = tmp395;
        assign tmp20 = mem_1[b3_w3];
        assign tmp432 = mem_3[tmp334];
    assign tmp40 = {shifted_w7[16], shifted_w7[17], shifted_w7[18], shifted_w7[19], shifted_w7[20], shifted_w7[21], shifted_w7[22], shifted_w7[23]};
    assign a2_w11 = tmp60;
        assign tmp2800 = mem_3[tmp2680];
        assign tmp528 = mem_3[tmp342];
    assign tmp1812 = tmp1872;
    assign tmp2774 = tmp2770 ^ tmp2773;
        assign tmp1299 = mem_3[tmp1212];
    assign tmp30 = w0 ^ xor_w3;
    assign tmp179 = concat_w27 ^ substituted_w27;
        assign tmp1652 = mem_3[tmp1510];
    assign tmp1522 = tmp1615;
    assign tmp2694 = tmp2787;
        assign tmp1180 = mem_1[tmp1148];
    assign tmp1230 = tmp1334;
    assign tmp1883 = tmp1879 ^ tmp1882;
    assign tmp1220 = {temp_14[16], temp_14[17], temp_14[18], temp_14[19], temp_14[20], temp_14[21], temp_14[22], temp_14[23]};
    assign temp_35 = tmp2896;
        assign tmp773 = mem_3[tmp631];
    assign tmp636 = {temp_6[0], temp_6[1], temp_6[2], temp_6[3], temp_6[4], temp_6[5], temp_6[6], temp_6[7]};
    assign tmp649 = tmp808;
    assign tmp2099 = {temp_26[16], temp_26[17], temp_26[18], temp_26[19], temp_26[20], temp_26[21], temp_26[22], temp_26[23]};
    assign tmp2775 = {tmp2774[0], tmp2774[1], tmp2774[2], tmp2774[3], tmp2774[4], tmp2774[5], tmp2774[6], tmp2774[7]};
    assign tmp539 = {tmp538[0], tmp538[1], tmp538[2], tmp538[3], tmp538[4], tmp538[5], tmp538[6], tmp538[7]};
    assign a3_w35 = tmp211;
    assign tmp1733 = {temp_20[72], temp_20[73], temp_20[74], temp_20[75], temp_20[76], temp_20[77], temp_20[78], temp_20[79]};
    assign tmp86 = {tmp83[8], tmp83[9], tmp83[10], tmp83[11], tmp83[12], tmp83[13], tmp83[14], tmp83[15]};
        assign tmp2640 = mem_1[tmp2608];
    assign tmp2072 = {temp_25[96], temp_25[97], temp_25[98], temp_25[99], temp_25[100], temp_25[101], temp_25[102], temp_25[103]};
    assign tmp2046 = tmp2062;
    assign tmp575 = tmp591;
        assign tmp2777 = mem_4[tmp2679];
    assign rc1_w27 = tmp174;
    assign tmp2235 = {tmp2234, tmp2094};
    assign tmp88 = {a2_w15, a3_w15, a4_w15, a1_w15};
    assign tmp112 = {tmp108[0], tmp108[1], tmp108[2], tmp108[3], tmp108[4], tmp108[5], tmp108[6], tmp108[7]};
    assign tmp2371 = {temp_29[48], temp_29[49], temp_29[50], temp_29[51], temp_29[52], temp_29[53], temp_29[54], temp_29[55]};
    assign tmp2560 = {tmp2559, tmp2393};
    assign tmp1503 = {temp_18[96], temp_18[97], temp_18[98], temp_18[99], temp_18[100], temp_18[101], temp_18[102], temp_18[103]};
    assign tmp1325 = tmp1323 ^ tmp1324;
    assign tmp1560 = {const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0, const1559_0};
    assign tmp2336 = tmp2352;
    assign tmp661 = {const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0, const660_0};
    assign tmp310 = {tmp278, tmp279, tmp280, tmp281, tmp282, tmp283, tmp284, tmp285, tmp286, tmp287, tmp288, tmp289, tmp290, tmp291, tmp292, tmp293};
    assign tmp1625 = {tmp1624, tmp1506};
    assign tmp1217 = {temp_14[40], temp_14[41], temp_14[42], temp_14[43], temp_14[44], temp_14[45], temp_14[46], temp_14[47]};
    assign tmp442 = tmp438 ^ tmp441;
    assign tmp955 = {tmp954, tmp917};
    assign tmp2244 = tmp2240 ^ tmp2243;
    assign tmp867 = tmp883;
        assign tmp1178 = mem_1[tmp1146];
    assign tmp735 = tmp731 ^ tmp734;
    assign tmp2258 = {const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0, const2257_0};
    assign tmp1317 = tmp1313 ^ tmp1316;
    assign tmp2488 = {tmp2487, tmp2383};
    assign xor_w3 = tmp29;
    assign tmp2838 = tmp2836 ^ tmp2837;
    assign tmp467 = {tmp466[0], tmp466[1], tmp466[2], tmp466[3], tmp466[4], tmp466[5], tmp466[6], tmp466[7]};
    assign input_wire_4 = temp_11;
    assign tmp1119 = {tmp1118, tmp926};
    assign tmp1778 = {temp_21[104], temp_21[105], temp_21[106], temp_21[107], temp_21[108], temp_21[109], temp_21[110], temp_21[111]};
    assign tmp2865 = {tmp2864, tmp2687};
    assign tmp686 = {tmp685, tmp622};
    assign tmp1116 = tmp1114 ^ tmp1115;
    assign tmp477 = {tmp476, tmp336};
    assign tmp1387 = {const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0, const1386_0};
    assign tmp285 = tmp301;
    assign tmp2361 = {tmp2329, tmp2330, tmp2331, tmp2332, tmp2333, tmp2334, tmp2335, tmp2336, tmp2337, tmp2338, tmp2339, tmp2340, tmp2341, tmp2342, tmp2343, tmp2344};
        assign tmp2166 = mem_3[tmp2090];
    assign tmp1953 = {const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0, const1952_0};
        assign tmp199 = mem_2[const198_8];
    assign tmp1929 = {const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0, const1928_0};
    assign tmp1732 = {temp_20[80], temp_20[81], temp_20[82], temp_20[83], temp_20[84], temp_20[85], temp_20[86], temp_20[87]};
        assign tmp1264 = mem_4[tmp1210];
        assign tmp2936 = mem_1[tmp2904];
    assign tmp635 = {temp_6[8], temp_6[9], temp_6[10], temp_6[11], temp_6[12], temp_6[13], temp_6[14], temp_6[15]};
        assign tmp1263 = mem_3[tmp1209];
    assign tmp161 = {tmp158[8], tmp158[9], tmp158[10], tmp158[11], tmp158[12], tmp158[13], tmp158[14], tmp158[15]};
    assign c4_w7 = tmp46;
    assign tmp291 = tmp307;
    assign tmp2198 = {const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0, const2197_0};
    assign tmp805 = {const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0, const804_0};
    assign tmp2700 = tmp2859;
    assign tmp1887 = tmp1885 ^ tmp1886;
    assign tmp2037 = tmp2053;
    assign tmp1111 = {tmp1110, tmp926};
    assign tmp1865 = {const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0, const1864_0};
        assign tmp118 = mem_1[b1_w19];
    assign tmp2665 = {temp_33[40], temp_33[41], temp_33[42], temp_33[43], temp_33[44], temp_33[45], temp_33[46], temp_33[47]};
    assign tmp1289 = tmp1287 ^ tmp1288;
    assign input_wire_2 = temp_3;
    assign tmp1565 = {tmp1564, tmp1501};
    assign tmp1458 = tmp1474;
    assign rc1_w11 = tmp74;
    assign tmp2760 = {const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0, const2759_0};
    assign tmp1088 = tmp1084 ^ tmp1087;
    assign temp_3 = tmp552;
    assign tmp2183 = {tmp2182, tmp2093};
        assign tmp445 = mem_4[tmp332];
    assign tmp215 = {shifted_w35[16], shifted_w35[17], shifted_w35[18], shifted_w35[19], shifted_w35[20], shifted_w35[21], shifted_w35[22], shifted_w35[23]};
    assign tmp210 = {tmp208[16], tmp208[17], tmp208[18], tmp208[19], tmp208[20], tmp208[21], tmp208[22], tmp208[23]};
    assign temp_18 = tmp1499;
    assign tmp231 = tmp230 ^ tmp206;
    assign tmp670 = {tmp669, tmp624};
    assign tmp1488 = {temp_17[80], temp_17[81], temp_17[82], temp_17[83], temp_17[84], temp_17[85], temp_17[86], temp_17[87]};
    assign tmp2144 = tmp2142 ^ tmp2143;
    assign tmp2175 = {tmp2174, tmp2093};
        assign tmp2358 = mem_1[tmp2326];
    assign tmp2172 = tmp2168 ^ tmp2171;
    assign tmp2030 = {temp_24[40], temp_24[41], temp_24[42], temp_24[43], temp_24[44], temp_24[45], temp_24[46], temp_24[47]};
    assign tmp695 = tmp691 ^ tmp694;
    assign tmp1221 = {temp_14[8], temp_14[9], temp_14[10], temp_14[11], temp_14[12], temp_14[13], temp_14[14], temp_14[15]};
    assign tmp1775 = {tmp1743, tmp1744, tmp1745, tmp1746, tmp1747, tmp1748, tmp1749, tmp1750, tmp1751, tmp1752, tmp1753, tmp1754, tmp1755, tmp1756, tmp1757, tmp1758};
    assign tmp1839 = tmp1837 ^ tmp1838;
        assign tmp1239 = mem_3[tmp1207];
        assign tmp2941 = mem_1[tmp2909];
    assign b2_w15 = tmp90;
        assign tmp2945 = mem_1[tmp2913];
    assign tmp1130 = {const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0, const1129_0};
    assign tmp1528 = tmp1687;
    assign tmp652 = tmp844;
    assign tmp2231 = {tmp2230, tmp2097};
    assign tmp1518 = tmp1567;
    assign tmp1248 = {tmp1247, tmp1210};
    assign tmp2603 = {tmp2395, tmp2396, tmp2397, tmp2398, tmp2399, tmp2400, tmp2401, tmp2402, tmp2403, tmp2404, tmp2405, tmp2406, tmp2407, tmp2408, tmp2409, tmp2410};
    assign tmp1685 = {tmp1684, tmp1515};
    assign tmp2127 = {tmp2126, tmp2089};
    assign tmp2491 = {const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0, const2490_0};
    assign tmp2109 = tmp2213;
    assign tmp10 = {w3[16], w3[17], w3[18], w3[19], w3[20], w3[21], w3[22], w3[23]};
    assign tmp1401 = tmp1397 ^ tmp1400;
    assign tmp2618 = {temp_32[24], temp_32[25], temp_32[26], temp_32[27], temp_32[28], temp_32[29], temp_32[30], temp_32[31]};
    assign shifted_w15 = tmp88;
        assign tmp1825 = mem_3[tmp1793];
    assign tmp1170 = tmp1186;
    assign tmp2095 = {temp_26[48], temp_26[49], temp_26[50], temp_26[51], temp_26[52], temp_26[53], temp_26[54], temp_26[55]};
    assign tmp2112 = tmp2249;
        assign tmp2812 = mem_3[tmp2681];
    assign a4_w39 = tmp237;
    assign tmp441 = {tmp440, tmp333};
    assign tmp632 = {temp_6[32], temp_6[33], temp_6[34], temp_6[35], temp_6[36], temp_6[37], temp_6[38], temp_6[39]};
    assign tmp1226 = tmp1286;
        assign tmp2645 = mem_1[tmp2613];
    assign tmp132 = tmp131 ^ tmp107;
    assign tmp1708 = {const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0, const1707_0};
    assign tmp1361 = tmp1359 ^ tmp1360;
    assign tmp1421 = tmp1419 ^ tmp1420;
    assign tmp920 = {temp_10[72], temp_10[73], temp_10[74], temp_10[75], temp_10[76], temp_10[77], temp_10[78], temp_10[79]};
    assign tmp1871 = tmp1867 ^ tmp1870;
    assign tmp2468 = {tmp2467, tmp2386};
    assign tmp1298 = {tmp1297[0], tmp1297[1], tmp1297[2], tmp1297[3], tmp1297[4], tmp1297[5], tmp1297[6], tmp1297[7]};
    assign tmp1056 = tmp1054 ^ tmp1055;
    assign tmp267 = {new_state[80], new_state[81], new_state[82], new_state[83], new_state[84], new_state[85], new_state[86], new_state[87]};
    assign tmp1040 = tmp1036 ^ tmp1039;
    assign tmp460 = {const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0, const459_0};
    assign tmp2609 = {temp_32[96], temp_32[97], temp_32[98], temp_32[99], temp_32[100], temp_32[101], temp_32[102], temp_32[103]};
        assign tmp1826 = mem_4[tmp1794];
        assign tmp493 = mem_4[tmp336];
        assign tmp2579 = mem_3[tmp2393];
    assign tmp2924 = tmp2940;
    assign tmp12 = {w3[0], w3[1], w3[2], w3[3], w3[4], w3[5], w3[6], w3[7]};
        assign tmp2055 = mem_1[tmp2023];
    assign tmp1155 = {temp_12[8], temp_12[9], temp_12[10], temp_12[11], temp_12[12], temp_12[13], temp_12[14], temp_12[15]};
    assign tmp2390 = {temp_30[32], temp_30[33], temp_30[34], temp_30[35], temp_30[36], temp_30[37], temp_30[38], temp_30[39]};
    assign tmp2840 = {const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0, const2839_0};
    assign tmp2464 = {tmp2463, tmp2385};
    assign tmp2691 = tmp2751;
        assign tmp599 = mem_1[tmp567];
    assign tmp1223 = tmp1250;
        assign tmp1383 = mem_3[tmp1219];
        assign tmp1921 = mem_3[tmp1801];
    assign c1_w35 = tmp218;
    assign tmp377 = {tmp376, tmp331};
    assign tmp2429 = tmp2425 ^ tmp2428;
    assign tmp669 = {const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0, const668_0};
    assign tmp847 = temp_7 ^ tmp846;
    assign tmp269 = {new_state[64], new_state[65], new_state[66], new_state[67], new_state[68], new_state[69], new_state[70], new_state[71]};
        assign tmp71 = mem_1[b4_w11];
    assign tmp1433 = temp_15 ^ tmp1432;
    assign tmp1614 = tmp1610 ^ tmp1613;
    assign tmp2071 = {temp_25[104], temp_25[105], temp_25[106], temp_25[107], temp_25[108], temp_25[109], temp_25[110], temp_25[111]};
    assign tmp2330 = tmp2346;
        assign tmp895 = mem_1[tmp863];
    assign tmp1896 = {tmp1895[0], tmp1895[1], tmp1895[2], tmp1895[3], tmp1895[4], tmp1895[5], tmp1895[6], tmp1895[7]};
    assign tmp213 = {a2_w35, a3_w35, a4_w35, a1_w35};
    assign tmp2658 = {temp_33[96], temp_33[97], temp_33[98], temp_33[99], temp_33[100], temp_33[101], temp_33[102], temp_33[103]};
    assign rc4_w39 = const252_0;
    assign tmp1520 = tmp1591;
    assign tmp1696 = {const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0, const1695_0};
    assign tmp763 = tmp761 ^ tmp762;
    assign tmp1842 = {tmp1841, tmp1796};
    assign tmp2040 = tmp2056;
    assign tmp503 = {tmp502[0], tmp502[1], tmp502[2], tmp502[3], tmp502[4], tmp502[5], tmp502[6], tmp502[7]};
    assign tmp1690 = tmp1688 ^ tmp1689;
    assign temp_39 = new_11;
    assign tmp1039 = {tmp1038, tmp920};
    assign tmp972 = tmp970 ^ tmp971;
    assign tmp1848 = {tmp1847[0], tmp1847[1], tmp1847[2], tmp1847[3], tmp1847[4], tmp1847[5], tmp1847[6], tmp1847[7]};
    assign tmp128 = {rc1_w19, rc2_w19, rc3_w19, rc4_w19};
    assign tmp1152 = {temp_12[32], temp_12[33], temp_12[34], temp_12[35], temp_12[36], temp_12[37], temp_12[38], temp_12[39]};
    assign tmp2019 = temp_23 ^ tmp2018;
    assign tmp1835 = tmp1831 ^ tmp1834;
    assign b3_w19 = tmp116;
    assign tmp1392 = {tmp1391, tmp1222};
    assign tmp268 = {new_state[72], new_state[73], new_state[74], new_state[75], new_state[76], new_state[77], new_state[78], new_state[79]};
        assign tmp1031 = mem_4[tmp918];
    assign tmp105 = tmp80 ^ xor_w15;
    assign tmp1949 = {const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0, const1948_0};
    assign temp_28 = new_8;
    assign tmp1915 = tmp1911 ^ tmp1914;
    assign tmp990 = {const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0, const989_0};
    assign tmp697 = {const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0, const696_0};
    assign tmp2912 = {temp_36[16], temp_36[17], temp_36[18], temp_36[19], temp_36[20], temp_36[21], temp_36[22], temp_36[23]};
        assign tmp305 = mem_1[tmp273];
    assign tmp1463 = tmp1479;
    assign tmp1755 = tmp1771;
    assign tmp117 = {shifted_w19[0], shifted_w19[1], shifted_w19[2], shifted_w19[3], shifted_w19[4], shifted_w19[5], shifted_w19[6], shifted_w19[7]};
    assign a4_w3 = tmp12;
    assign tmp2405 = tmp2542;
    assign tmp1399 = {const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0, const1398_0};
    assign tmp879 = tmp895;
    assign c1_w11 = tmp68;
    assign tmp719 = tmp715 ^ tmp718;
        assign tmp1114 = mem_3[tmp928];
    assign shifted_w7 = tmp38;
    assign tmp41 = {shifted_w7[8], shifted_w7[9], shifted_w7[10], shifted_w7[11], shifted_w7[12], shifted_w7[13], shifted_w7[14], shifted_w7[15]};
    assign tmp1515 = {temp_18[0], temp_18[1], temp_18[2], temp_18[3], temp_18[4], temp_18[5], temp_18[6], temp_18[7]};
    assign tmp2278 = {const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0, const2277_0};
    assign tmp2425 = tmp2423 ^ tmp2424;
        assign tmp2861 = mem_4[tmp2686];
    assign tmp2572 = {tmp2571, tmp2394};
        assign tmp1592 = mem_3[tmp1505];
    assign tmp1973 = {const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0, const1972_0};
    assign tmp771 = tmp767 ^ tmp770;
    assign tmp1536 = {const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0, const1535_0};
    assign tmp2620 = {temp_32[8], temp_32[9], temp_32[10], temp_32[11], temp_32[12], temp_32[13], temp_32[14], temp_32[15]};
    assign tmp2276 = tmp2274 ^ tmp2275;
    assign tmp904 = {temp_9[64], temp_9[65], temp_9[66], temp_9[67], temp_9[68], temp_9[69], temp_9[70], temp_9[71]};
        assign tmp738 = mem_4[tmp625];
    assign tmp829 = {const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0, const828_0};
    assign tmp486 = tmp482 ^ tmp485;
    assign tmp2533 = tmp2531 ^ tmp2532;
    assign tmp2207 = {tmp2206, tmp2091};
    assign tmp2136 = tmp2132 ^ tmp2135;
    assign tmp2561 = tmp2557 ^ tmp2560;
    assign tmp2712 = {const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0, const2711_0};
    assign b3_w3 = tmp16;
    assign tmp2445 = tmp2441 ^ tmp2444;
    assign tmp276 = {new_state[8], new_state[9], new_state[10], new_state[11], new_state[12], new_state[13], new_state[14], new_state[15]};
    assign c2_w35 = tmp219;
    assign tmp619 = {temp_5[0], temp_5[1], temp_5[2], temp_5[3], temp_5[4], temp_5[5], temp_5[6], temp_5[7]};
    assign tmp1296 = {tmp1295, tmp1214};
        assign tmp1184 = mem_1[tmp1152];
    assign tmp870 = tmp886;
    assign tmp2957 = {temp_37[48], temp_37[49], temp_37[50], temp_37[51], temp_37[52], temp_37[53], temp_37[54], temp_37[55]};
    assign b2_w11 = tmp65;
        assign tmp2226 = mem_3[tmp2095];
    assign tmp7 = {aes_key[32], aes_key[33], aes_key[34], aes_key[35], aes_key[36], aes_key[37], aes_key[38], aes_key[39], aes_key[40], aes_key[41], aes_key[42], aes_key[43], aes_key[44], aes_key[45], aes_key[46], aes_key[47], aes_key[48], aes_key[49], aes_key[50], aes_key[51], aes_key[52], aes_key[53], aes_key[54], aes_key[55], aes_key[56], aes_key[57], aes_key[58], aes_key[59], aes_key[60], aes_key[61], aes_key[62], aes_key[63]};
    assign tmp1238 = tmp1430;
    assign tmp2291 = {tmp2290, tmp2098};
        assign tmp1762 = mem_1[tmp1730];
    assign tmp2587 = {const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0, const2586_0};
    assign tmp340 = {temp_2[24], temp_2[25], temp_2[26], temp_2[27], temp_2[28], temp_2[29], temp_2[30], temp_2[31]};
    assign tmp2148 = tmp2144 ^ tmp2147;
    assign tmp368 = {const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0, const367_0};
    assign tmp747 = tmp743 ^ tmp746;
    assign tmp1292 = {tmp1291, tmp1213};
    assign tmp2069 = {temp_25[120], temp_25[121], temp_25[122], temp_25[123], temp_25[124], temp_25[125], temp_25[126], temp_25[127]};
    assign tmp578 = tmp594;
    assign tmp766 = {tmp765, tmp632};
    assign tmp1827 = tmp1825 ^ tmp1826;
    assign tmp753 = {const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0, const752_0};
    assign tmp1983 = tmp1981 ^ tmp1982;
    assign tmp335 = {temp_2[64], temp_2[65], temp_2[66], temp_2[67], temp_2[68], temp_2[69], temp_2[70], temp_2[71]};
    assign tmp2259 = {tmp2258, tmp2096};
        assign tmp1176 = mem_1[tmp1144];
    assign tmp1821 = tmp1980;
    assign tmp2024 = {temp_24[88], temp_24[89], temp_24[90], temp_24[91], temp_24[92], temp_24[93], temp_24[94], temp_24[95]};
    assign tmp318 = {temp_1[64], temp_1[65], temp_1[66], temp_1[67], temp_1[68], temp_1[69], temp_1[70], temp_1[71]};
    assign tmp205 = tmp180 ^ xor_w31;
    assign tmp2697 = tmp2823;
    assign tmp2876 = {const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0, const2875_0};
    assign tmp2026 = {temp_24[72], temp_24[73], temp_24[74], temp_24[75], temp_24[76], temp_24[77], temp_24[78], temp_24[79]};
    assign tmp2007 = tmp2005 ^ tmp2006;
    assign tmp1543 = {tmp1542[0], tmp1542[1], tmp1542[2], tmp1542[3], tmp1542[4], tmp1542[5], tmp1542[6], tmp1542[7]};
    assign c2_w19 = tmp119;
    assign tmp2138 = {const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0, const2137_0};
        assign tmp2349 = mem_1[tmp2317];
    assign tmp2754 = tmp2752 ^ tmp2753;
    assign tmp1875 = tmp1873 ^ tmp1874;
        assign tmp2178 = mem_3[tmp2091];
    assign tmp609 = {temp_5[80], temp_5[81], temp_5[82], temp_5[83], temp_5[84], temp_5[85], temp_5[86], temp_5[87]};
    assign tmp2784 = {const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0, const2783_0};
    assign tmp2273 = {tmp2272[0], tmp2272[1], tmp2272[2], tmp2272[3], tmp2272[4], tmp2272[5], tmp2272[6], tmp2272[7]};
    assign tmp501 = {tmp500, tmp338};
    assign tmp2085 = {tmp2069, tmp2074, tmp2079, tmp2084, tmp2073, tmp2078, tmp2083, tmp2072, tmp2077, tmp2082, tmp2071, tmp2076, tmp2081, tmp2070, tmp2075, tmp2080};
    assign tmp1261 = tmp1257 ^ tmp1260;
    assign tmp794 = {tmp793, tmp631};
    assign tmp1351 = {const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0, const1350_0};
    assign tmp351 = tmp455;
    assign tmp2613 = {temp_32[64], temp_32[65], temp_32[66], temp_32[67], temp_32[68], temp_32[69], temp_32[70], temp_32[71]};
    assign tmp992 = tmp988 ^ tmp991;
        assign tmp2484 = mem_4[tmp2386];
    assign tmp1702 = tmp1700 ^ tmp1701;
    assign tmp1660 = {const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0, const1659_0};
    assign tmp165 = {shifted_w27[16], shifted_w27[17], shifted_w27[18], shifted_w27[19], shifted_w27[20], shifted_w27[21], shifted_w27[22], shifted_w27[23]};
    assign tmp473 = {tmp472, tmp339};
    assign tmp2828 = {const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0, const2827_0};
    assign tmp639 = tmp688;
    assign tmp2313 = {temp_28[120], temp_28[121], temp_28[122], temp_28[123], temp_28[124], temp_28[125], temp_28[126], temp_28[127]};
    assign tmp1100 = tmp1096 ^ tmp1099;
    assign tmp60 = {tmp58[16], tmp58[17], tmp58[18], tmp58[19], tmp58[20], tmp58[21], tmp58[22], tmp58[23]};
    assign b1_w35 = tmp214;
    assign tmp1845 = {const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0, const1844_0};
    assign tmp2362 = {temp_29[120], temp_29[121], temp_29[122], temp_29[123], temp_29[124], temp_29[125], temp_29[126], temp_29[127]};
    assign tmp2617 = {temp_32[32], temp_32[33], temp_32[34], temp_32[35], temp_32[36], temp_32[37], temp_32[38], temp_32[39]};
    assign tmp793 = {const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0, const792_0};
    assign tmp378 = tmp374 ^ tmp377;
    assign tmp1328 = {tmp1327, tmp1212};
    assign temp_24 = new_7;
    assign tmp1661 = {tmp1660, tmp1509};
    assign tmp79 = concat_w11 ^ substituted_w11;
        assign tmp1419 = mem_3[tmp1222];
    assign tmp334 = {temp_2[72], temp_2[73], temp_2[74], temp_2[75], temp_2[76], temp_2[77], temp_2[78], temp_2[79]};
    assign tmp1285 = tmp1281 ^ tmp1284;
    assign tmp2566 = {tmp2565[0], tmp2565[1], tmp2565[2], tmp2565[3], tmp2565[4], tmp2565[5], tmp2565[6], tmp2565[7]};
    assign rc4_w15 = const102_0;
    assign tmp97 = {c1_w15, c2_w15, c3_w15, c4_w15};
    assign tmp1941 = {const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0, const1940_0};
    assign tmp116 = {shifted_w19[8], shifted_w19[9], shifted_w19[10], shifted_w19[11], shifted_w19[12], shifted_w19[13], shifted_w19[14], shifted_w19[15]};
    assign tmp2730 = tmp2728 ^ tmp2729;
    assign tmp184 = {tmp183[24], tmp183[25], tmp183[26], tmp183[27], tmp183[28], tmp183[29], tmp183[30], tmp183[31]};
    assign tmp1521 = tmp1603;
    assign tmp417 = {tmp416, tmp335};
    assign tmp1343 = {const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0, const1342_0};
    assign tmp743 = tmp739 ^ tmp742;
    assign tmp1682 = tmp1678 ^ tmp1681;
    assign tmp858 = {temp_8[40], temp_8[41], temp_8[42], temp_8[43], temp_8[44], temp_8[45], temp_8[46], temp_8[47]};
    assign concat_w35 = tmp228;
    assign tmp2792 = {const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0, const2791_0};
    assign tmp2772 = {const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0, const2771_0};
        assign tmp1933 = mem_3[tmp1802];
    assign tmp923 = {temp_10[48], temp_10[49], temp_10[50], temp_10[51], temp_10[52], temp_10[53], temp_10[54], temp_10[55]};
    assign tmp815 = tmp811 ^ tmp814;
    assign tmp914 = {temp_10[120], temp_10[121], temp_10[122], temp_10[123], temp_10[124], temp_10[125], temp_10[126], temp_10[127]};
    assign tmp1034 = {const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0, const1033_0};
    assign tmp868 = tmp884;
        assign tmp809 = mem_3[tmp634];
    assign tmp2180 = tmp2178 ^ tmp2179;
    assign tmp1817 = tmp1932;
        assign tmp146 = mem_1[b4_w23];
    assign tmp2373 = {temp_29[32], temp_29[33], temp_29[34], temp_29[35], temp_29[36], temp_29[37], temp_29[38], temp_29[39]};
    assign b1_w19 = tmp114;
    assign tmp1724 = {tmp1516, tmp1517, tmp1518, tmp1519, tmp1520, tmp1521, tmp1522, tmp1523, tmp1524, tmp1525, tmp1526, tmp1527, tmp1528, tmp1529, tmp1530, tmp1531};
    assign tmp2383 = {temp_30[88], temp_30[89], temp_30[90], temp_30[91], temp_30[92], temp_30[93], temp_30[94], temp_30[95]};
    assign w6 = tmp32;
    assign rc1_w31 = tmp199;
    assign tmp2571 = {const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0, const2570_0};
    assign tmp1243 = {const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0, const1242_0};
    assign tmp1748 = tmp1764;
    assign tmp1600 = {const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0, const1599_0};
    assign tmp2113 = tmp2261;
        assign tmp714 = mem_4[tmp627];
    assign tmp1483 = {temp_17[120], temp_17[121], temp_17[122], temp_17[123], temp_17[124], temp_17[125], temp_17[126], temp_17[127]};
    assign tmp715 = tmp713 ^ tmp714;
    assign tmp1603 = {tmp1602[0], tmp1602[1], tmp1602[2], tmp1602[3], tmp1602[4], tmp1602[5], tmp1602[6], tmp1602[7]};
    assign temp_38 = tmp2964;
    assign tmp1944 = {tmp1943[0], tmp1943[1], tmp1943[2], tmp1943[3], tmp1943[4], tmp1943[5], tmp1943[6], tmp1943[7]};
    assign tmp2679 = {temp_34[64], temp_34[65], temp_34[66], temp_34[67], temp_34[68], temp_34[69], temp_34[70], temp_34[71]};
    assign rc1_w19 = tmp124;
    assign tmp1833 = {const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0, const1832_0};
        assign tmp295 = mem_1[tmp263];
    assign tmp683 = tmp679 ^ tmp682;
    assign tmp754 = {tmp753, tmp631};
    assign tmp450 = tmp446 ^ tmp449;
    assign tmp2569 = tmp2567 ^ tmp2568;
    assign tmp187 = {tmp183[0], tmp183[1], tmp183[2], tmp183[3], tmp183[4], tmp183[5], tmp183[6], tmp183[7]};
    assign tmp1413 = tmp1409 ^ tmp1412;
        assign tmp246 = mem_1[b4_w39];
    assign concat_w15 = tmp103;
    assign a3_w7 = tmp36;
    assign tmp2565 = tmp2561 ^ tmp2564;
    assign tmp1648 = {const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0, const1647_0};
    assign tmp1457 = tmp1473;
    assign tmp114 = {shifted_w19[24], shifted_w19[25], shifted_w19[26], shifted_w19[27], shifted_w19[28], shifted_w19[29], shifted_w19[30], shifted_w19[31]};
        assign tmp18 = mem_1[b1_w3];
    assign tmp901 = {temp_9[88], temp_9[89], temp_9[90], temp_9[91], temp_9[92], temp_9[93], temp_9[94], temp_9[95]};
    assign tmp604 = {temp_5[120], temp_5[121], temp_5[122], temp_5[123], temp_5[124], temp_5[125], temp_5[126], temp_5[127]};
    assign tmp1495 = {temp_17[24], temp_17[25], temp_17[26], temp_17[27], temp_17[28], temp_17[29], temp_17[30], temp_17[31]};
    assign tmp2378 = {tmp2362, tmp2367, tmp2372, tmp2377, tmp2366, tmp2371, tmp2376, tmp2365, tmp2370, tmp2375, tmp2364, tmp2369, tmp2374, tmp2363, tmp2368, tmp2373};
    assign tmp1236 = tmp1406;
    assign tmp2135 = {tmp2134, tmp2089};
    assign tmp2015 = tmp2011 ^ tmp2014;
    assign tmp1277 = tmp1275 ^ tmp1276;
    assign tmp2098 = {temp_26[24], temp_26[25], temp_26[26], temp_26[27], temp_26[28], temp_26[29], temp_26[30], temp_26[31]};
    assign tmp1005 = {tmp1004[0], tmp1004[1], tmp1004[2], tmp1004[3], tmp1004[4], tmp1004[5], tmp1004[6], tmp1004[7]};
    assign b4_w39 = tmp242;
        assign tmp1568 = mem_3[tmp1503];
    assign tmp139 = {shifted_w23[24], shifted_w23[25], shifted_w23[26], shifted_w23[27], shifted_w23[28], shifted_w23[29], shifted_w23[30], shifted_w23[31]};
    assign tmp2674 = {temp_34[104], temp_34[105], temp_34[106], temp_34[107], temp_34[108], temp_34[109], temp_34[110], temp_34[111]};
    assign tmp2212 = tmp2208 ^ tmp2211;
    assign tmp906 = {temp_9[48], temp_9[49], temp_9[50], temp_9[51], temp_9[52], temp_9[53], temp_9[54], temp_9[55]};
    assign tmp564 = {temp_4[48], temp_4[49], temp_4[50], temp_4[51], temp_4[52], temp_4[53], temp_4[54], temp_4[55]};
        assign tmp1664 = mem_3[tmp1511];
    assign tmp618 = {temp_5[8], temp_5[9], temp_5[10], temp_5[11], temp_5[12], temp_5[13], temp_5[14], temp_5[15]};
    assign tmp1260 = {tmp1259, tmp1207};
    assign b1_w39 = tmp239;
        assign tmp2006 = mem_4[tmp1805];
        assign tmp1773 = mem_1[tmp1741];
    assign tmp2338 = tmp2354;
        assign tmp218 = mem_1[b1_w35];
    assign tmp1189 = {tmp1157, tmp1158, tmp1159, tmp1160, tmp1161, tmp1162, tmp1163, tmp1164, tmp1165, tmp1166, tmp1167, tmp1168, tmp1169, tmp1170, tmp1171, tmp1172};
        assign tmp1763 = mem_1[tmp1731];
    assign tmp855 = {temp_8[64], temp_8[65], temp_8[66], temp_8[67], temp_8[68], temp_8[69], temp_8[70], temp_8[71]};
    assign tmp2473 = tmp2471 ^ tmp2472;
    assign tmp2874 = tmp2872 ^ tmp2873;
        assign tmp1759 = mem_1[tmp1727];
    assign new_6 = tmp1726;
    assign tmp2616 = {temp_32[40], temp_32[41], temp_32[42], temp_32[43], temp_32[44], temp_32[45], temp_32[46], temp_32[47]};
        assign tmp2939 = mem_1[tmp2907];
    assign tmp784 = {tmp783[0], tmp783[1], tmp783[2], tmp783[3], tmp783[4], tmp783[5], tmp783[6], tmp783[7]};
    assign tmp2751 = {tmp2750[0], tmp2750[1], tmp2750[2], tmp2750[3], tmp2750[4], tmp2750[5], tmp2750[6], tmp2750[7]};
    assign tmp1253 = tmp1251 ^ tmp1252;
    assign tmp2094 = {temp_26[56], temp_26[57], temp_26[58], temp_26[59], temp_26[60], temp_26[61], temp_26[62], temp_26[63]};
    assign tmp2045 = tmp2061;
    assign tmp2151 = {tmp2150, tmp2087};
        assign tmp1177 = mem_1[tmp1145];
    assign c4_w15 = tmp96;
    assign tmp623 = {temp_6[104], temp_6[105], temp_6[106], temp_6[107], temp_6[108], temp_6[109], temp_6[110], temp_6[111]};
    assign tmp717 = {const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0, const716_0};
    assign b2_w39 = tmp240;
    assign tmp2117 = tmp2309;
    assign c3_w31 = tmp195;
    assign tmp745 = {const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0, const744_0};
    assign tmp999 = {tmp998, tmp920};
    assign tmp546 = tmp542 ^ tmp545;
    assign tmp2325 = {temp_28[24], temp_28[25], temp_28[26], temp_28[27], temp_28[28], temp_28[29], temp_28[30], temp_28[31]};
        assign tmp2544 = mem_4[tmp2387];
    assign tmp322 = {temp_1[32], temp_1[33], temp_1[34], temp_1[35], temp_1[36], temp_1[37], temp_1[38], temp_1[39]};
    assign tmp1224 = tmp1262;
    assign tmp1036 = tmp1032 ^ tmp1035;
    assign tmp1228 = tmp1310;
    assign tmp864 = tmp880;
    assign tmp2744 = {const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0, const2743_0};
    assign tmp1578 = tmp1574 ^ tmp1577;
    assign tmp1564 = {const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0, const1563_0};
        assign tmp2580 = mem_4[tmp2394];
    assign tmp2762 = tmp2758 ^ tmp2761;
    assign tmp1714 = tmp1712 ^ tmp1713;
    assign tmp1349 = tmp1347 ^ tmp1348;
    assign tmp9 = {w3[24], w3[25], w3[26], w3[27], w3[28], w3[29], w3[30], w3[31]};
        assign tmp2495 = mem_3[tmp2386];
    assign tmp2100 = {temp_26[8], temp_26[9], temp_26[10], temp_26[11], temp_26[12], temp_26[13], temp_26[14], temp_26[15]};
        assign tmp2641 = mem_1[tmp2609];
    assign tmp111 = {tmp108[8], tmp108[9], tmp108[10], tmp108[11], tmp108[12], tmp108[13], tmp108[14], tmp108[15]};
    assign tmp1297 = tmp1293 ^ tmp1296;
        assign tmp1396 = mem_4[tmp1221];
    assign a3_w31 = tmp186;
    assign tmp524 = {const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0, const523_0};
    assign tmp2947 = {tmp2915, tmp2916, tmp2917, tmp2918, tmp2919, tmp2920, tmp2921, tmp2922, tmp2923, tmp2924, tmp2925, tmp2926, tmp2927, tmp2928, tmp2929, tmp2930};
    assign tmp934 = tmp1005;
    assign tmp679 = tmp677 ^ tmp678;
    assign a1_w7 = tmp34;
        assign tmp421 = mem_4[tmp334];
    assign tmp1554 = tmp1550 ^ tmp1553;
    assign tmp1255 = {const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0, const1254_0};
    assign tmp2260 = tmp2256 ^ tmp2259;
    assign tmp331 = {temp_2[96], temp_2[97], temp_2[98], temp_2[99], temp_2[100], temp_2[101], temp_2[102], temp_2[103]};
    assign b3_w35 = tmp216;
        assign tmp1173 = mem_1[tmp1141];
        assign tmp456 = mem_3[tmp336];
    assign tmp2678 = {temp_34[72], temp_34[73], temp_34[74], temp_34[75], temp_34[76], temp_34[77], temp_34[78], temp_34[79]};
    assign tmp1032 = tmp1030 ^ tmp1031;
    assign tmp1060 = tmp1056 ^ tmp1059;
        assign tmp2813 = mem_4[tmp2682];
    assign a3_w11 = tmp61;
    assign tmp2031 = {temp_24[32], temp_24[33], temp_24[34], temp_24[35], temp_24[36], temp_24[37], temp_24[38], temp_24[39]};
    assign tmp727 = tmp725 ^ tmp726;
    assign tmp2959 = {temp_37[32], temp_37[33], temp_37[34], temp_37[35], temp_37[36], temp_37[37], temp_37[38], temp_37[39]};
    assign b3_w39 = tmp241;
        assign tmp1471 = mem_1[tmp1439];
    assign tmp1793 = {temp_22[120], temp_22[121], temp_22[122], temp_22[123], temp_22[124], temp_22[125], temp_22[126], temp_22[127]};
        assign tmp1653 = mem_4[tmp1511];
        assign tmp2062 = mem_1[tmp2030];
    assign tmp608 = {temp_5[88], temp_5[89], temp_5[90], temp_5[91], temp_5[92], temp_5[93], temp_5[94], temp_5[95]};
        assign tmp2262 = mem_3[tmp2098];
    assign tmp1608 = {const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0, const1607_0};
    assign tmp2333 = tmp2349;
    assign tmp2539 = {const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0, const2538_0};
    assign tmp2139 = {tmp2138, tmp2086};
    assign tmp1811 = tmp1860;
    assign tmp2469 = tmp2465 ^ tmp2468;
    assign tmp2799 = {tmp2798[0], tmp2798[1], tmp2798[2], tmp2798[3], tmp2798[4], tmp2798[5], tmp2798[6], tmp2798[7]};
    assign tmp693 = {const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0, const692_0};
    assign tmp2232 = tmp2228 ^ tmp2231;
    assign tmp664 = {tmp663[0], tmp663[1], tmp663[2], tmp663[3], tmp663[4], tmp663[5], tmp663[6], tmp663[7]};
    assign xor_w15 = tmp104;
    assign tmp2523 = {const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0, const2522_0};
        assign tmp505 = mem_4[tmp341];
    assign tmp2527 = {const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0, const2526_0};
    assign concat_w11 = tmp78;
    assign tmp630 = {temp_6[48], temp_6[49], temp_6[50], temp_6[51], temp_6[52], temp_6[53], temp_6[54], temp_6[55]};
    assign b4_w19 = tmp117;
        assign tmp2056 = mem_1[tmp2024];
    assign temp_17 = tmp1482;
    assign tmp533 = {tmp532, tmp340};
    assign tmp2595 = {const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0, const2594_0};
    assign tmp2340 = tmp2356;
    assign c4_w27 = tmp171;
        assign tmp1468 = mem_1[tmp1436];
    assign tmp648 = tmp796;
        assign tmp1874 = mem_4[tmp1798];
    assign tmp2184 = tmp2180 ^ tmp2183;
    assign tmp848 = {temp_8[120], temp_8[121], temp_8[122], temp_8[123], temp_8[124], temp_8[125], temp_8[126], temp_8[127]};
    assign rc4_w11 = const77_0;
    assign tmp1858 = {tmp1857, tmp1794};
    assign tmp2387 = {temp_30[56], temp_30[57], temp_30[58], temp_30[59], temp_30[60], temp_30[61], temp_30[62], temp_30[63]};
    assign c4_w3 = tmp21;
    assign rc3_w19 = const126_0;
    assign tmp262 = {new_state[120], new_state[121], new_state[122], new_state[123], new_state[124], new_state[125], new_state[126], new_state[127]};
        assign tmp1838 = mem_4[tmp1795];
    assign tmp162 = {tmp158[0], tmp158[1], tmp158[2], tmp158[3], tmp158[4], tmp158[5], tmp158[6], tmp158[7]};
    assign tmp2850 = tmp2848 ^ tmp2849;
    assign tmp2315 = {temp_28[104], temp_28[105], temp_28[106], temp_28[107], temp_28[108], temp_28[109], temp_28[110], temp_28[111]};
    assign tmp2830 = tmp2826 ^ tmp2829;
    assign tmp2219 = {tmp2218, tmp2096};
    assign tmp2479 = {const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0, const2478_0};
    assign tmp1122 = {const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0, const1121_0};
    assign tmp2398 = tmp2458;
    assign tmp2536 = {tmp2535, tmp2387};
    assign tmp1016 = tmp1012 ^ tmp1015;
    assign tmp1920 = {tmp1919[0], tmp1919[1], tmp1919[2], tmp1919[3], tmp1919[4], tmp1919[5], tmp1919[6], tmp1919[7]};
        assign tmp504 = mem_3[tmp340];
    assign tmp638 = tmp676;
    assign tmp412 = {const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0, const411_0};
        assign tmp2653 = mem_1[tmp2621];
    assign tmp2428 = {tmp2427, tmp2382};
    assign tmp1978 = {tmp1977, tmp1808};
    assign tmp1451 = tmp1467;
    assign tmp513 = {tmp512, tmp343};
    assign tmp214 = {shifted_w35[24], shifted_w35[25], shifted_w35[26], shifted_w35[27], shifted_w35[28], shifted_w35[29], shifted_w35[30], shifted_w35[31]};
    assign tmp1549 = {tmp1548, tmp1503};
    assign tmp2768 = {const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0, const2767_0};
        assign tmp46 = mem_1[b4_w7];
    assign tmp8 = {aes_key[0], aes_key[1], aes_key[2], aes_key[3], aes_key[4], aes_key[5], aes_key[6], aes_key[7], aes_key[8], aes_key[9], aes_key[10], aes_key[11], aes_key[12], aes_key[13], aes_key[14], aes_key[15], aes_key[16], aes_key[17], aes_key[18], aes_key[19], aes_key[20], aes_key[21], aes_key[22], aes_key[23], aes_key[24], aes_key[25], aes_key[26], aes_key[27], aes_key[28], aes_key[29], aes_key[30], aes_key[31]};
    assign tmp510 = tmp506 ^ tmp509;
    assign tmp941 = tmp1089;
    assign tmp2271 = {tmp2270, tmp2101};
        assign tmp1469 = mem_1[tmp1437];
    assign tmp2018 = {expanded_key[512], expanded_key[513], expanded_key[514], expanded_key[515], expanded_key[516], expanded_key[517], expanded_key[518], expanded_key[519], expanded_key[520], expanded_key[521], expanded_key[522], expanded_key[523], expanded_key[524], expanded_key[525], expanded_key[526], expanded_key[527], expanded_key[528], expanded_key[529], expanded_key[530], expanded_key[531], expanded_key[532], expanded_key[533], expanded_key[534], expanded_key[535], expanded_key[536], expanded_key[537], expanded_key[538], expanded_key[539], expanded_key[540], expanded_key[541], expanded_key[542], expanded_key[543], expanded_key[544], expanded_key[545], expanded_key[546], expanded_key[547], expanded_key[548], expanded_key[549], expanded_key[550], expanded_key[551], expanded_key[552], expanded_key[553], expanded_key[554], expanded_key[555], expanded_key[556], expanded_key[557], expanded_key[558], expanded_key[559], expanded_key[560], expanded_key[561], expanded_key[562], expanded_key[563], expanded_key[564], expanded_key[565], expanded_key[566], expanded_key[567], expanded_key[568], expanded_key[569], expanded_key[570], expanded_key[571], expanded_key[572], expanded_key[573], expanded_key[574], expanded_key[575], expanded_key[576], expanded_key[577], expanded_key[578], expanded_key[579], expanded_key[580], expanded_key[581], expanded_key[582], expanded_key[583], expanded_key[584], expanded_key[585], expanded_key[586], expanded_key[587], expanded_key[588], expanded_key[589], expanded_key[590], expanded_key[591], expanded_key[592], expanded_key[593], expanded_key[594], expanded_key[595], expanded_key[596], expanded_key[597], expanded_key[598], expanded_key[599], expanded_key[600], expanded_key[601], expanded_key[602], expanded_key[603], expanded_key[604], expanded_key[605], expanded_key[606], expanded_key[607], expanded_key[608], expanded_key[609], expanded_key[610], expanded_key[611], expanded_key[612], expanded_key[613], expanded_key[614], expanded_key[615], expanded_key[616], expanded_key[617], expanded_key[618], expanded_key[619], expanded_key[620], expanded_key[621], expanded_key[622], expanded_key[623], expanded_key[624], expanded_key[625], expanded_key[626], expanded_key[627], expanded_key[628], expanded_key[629], expanded_key[630], expanded_key[631], expanded_key[632], expanded_key[633], expanded_key[634], expanded_key[635], expanded_key[636], expanded_key[637], expanded_key[638], expanded_key[639]};
        assign tmp1765 = mem_1[tmp1733];
        assign tmp2179 = mem_4[tmp2092];
    assign tmp2366 = {temp_29[88], temp_29[89], temp_29[90], temp_29[91], temp_29[92], temp_29[93], temp_29[94], temp_29[95]};
        assign tmp588 = mem_1[tmp556];
    assign tmp1654 = tmp1652 ^ tmp1653;
    assign tmp2147 = {tmp2146, tmp2086};
    assign tmp676 = {tmp675[0], tmp675[1], tmp675[2], tmp675[3], tmp675[4], tmp675[5], tmp675[6], tmp675[7]};
    assign new_4 = tmp1140;
    assign tmp2384 = {temp_30[80], temp_30[81], temp_30[82], temp_30[83], temp_30[84], temp_30[85], temp_30[86], temp_30[87]};
    assign tmp527 = {tmp526[0], tmp526[1], tmp526[2], tmp526[3], tmp526[4], tmp526[5], tmp526[6], tmp526[7]};
    assign tmp837 = {const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0, const836_0};
    assign tmp2746 = tmp2742 ^ tmp2745;
    assign tmp66 = {shifted_w11[8], shifted_w11[9], shifted_w11[10], shifted_w11[11], shifted_w11[12], shifted_w11[13], shifted_w11[14], shifted_w11[15]};
    assign tmp2111 = tmp2237;
    assign tmp108 = tmp107 ^ tmp83;
    assign tmp2087 = {temp_26[112], temp_26[113], temp_26[114], temp_26[115], temp_26[116], temp_26[117], temp_26[118], temp_26[119]};
    assign a3_w23 = tmp136;
    assign tmp532 = {const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0, const531_0};
    assign tmp655 = tmp653 ^ tmp654;
    assign tmp924 = {temp_10[40], temp_10[41], temp_10[42], temp_10[43], temp_10[44], temp_10[45], temp_10[46], temp_10[47]};
    assign substituted_w11 = tmp72;
    assign tmp147 = {c1_w23, c2_w23, c3_w23, c4_w23};
    assign tmp781 = {const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0, const780_0};
    assign tmp1626 = tmp1622 ^ tmp1625;
    assign tmp2804 = {const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0, const2803_0};
    assign tmp2079 = {temp_25[40], temp_25[41], temp_25[42], temp_25[43], temp_25[44], temp_25[45], temp_25[46], temp_25[47]};
    assign tmp703 = tmp701 ^ tmp702;
    assign tmp2035 = {temp_24[0], temp_24[1], temp_24[2], temp_24[3], temp_24[4], temp_24[5], temp_24[6], temp_24[7]};
    assign rc4_w27 = const177_0;
    assign tmp2206 = {const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0, const2205_0};
    assign tmp1158 = tmp1174;
    assign tmp13 = {a2_w3, a3_w3, a4_w3, a1_w3};
    assign tmp2415 = {const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0, const2414_0};
        assign tmp2801 = mem_4[tmp2681];
    assign tmp259 = {w0, w1, w2, w3, w4, w5, w6, w7, tmp55, tmp56, tmp57, tmp58, tmp80, tmp81, tmp82, tmp83, tmp105, tmp106, tmp107, tmp108, tmp130, tmp131, tmp132, tmp133, tmp155, tmp156, tmp157, tmp158, tmp180, tmp181, tmp182, tmp183, tmp205, tmp206, tmp207, tmp208, tmp230, tmp231, tmp232, tmp233, tmp255, tmp256, tmp257, tmp258};
    assign tmp2380 = {temp_30[112], temp_30[113], temp_30[114], temp_30[115], temp_30[116], temp_30[117], temp_30[118], temp_30[119]};
    assign tmp1524 = tmp1639;
    assign tmp954 = {const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0, const953_0};
    assign c2_w11 = tmp69;
        assign tmp2143 = mem_4[tmp2089];
        assign tmp2872 = mem_3[tmp2686];
    assign tmp426 = tmp422 ^ tmp425;
    assign tmp940 = tmp1077;
    assign tmp2255 = {tmp2254, tmp2095};
    assign tmp364 = {const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0, const363_0};
    assign tmp739 = tmp737 ^ tmp738;
    assign tmp1492 = {temp_17[48], temp_17[49], temp_17[50], temp_17[51], temp_17[52], temp_17[53], temp_17[54], temp_17[55]};
        assign tmp2436 = mem_4[tmp2382];
    assign tmp1697 = {tmp1696, tmp1512};
        assign tmp45 = mem_1[b3_w7];
    assign tmp2042 = tmp2058;
    assign tmp2432 = {tmp2431, tmp2379};
    assign tmp2020 = {temp_24[120], temp_24[121], temp_24[122], temp_24[123], temp_24[124], temp_24[125], temp_24[126], temp_24[127]};
    assign tmp413 = {tmp412, tmp334};
    assign new_5 = tmp1433;
        assign tmp221 = mem_1[b4_w35];
    assign tmp520 = {const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0, const519_0};
    assign tmp1529 = tmp1699;
    assign tmp389 = {tmp388, tmp328};
        assign tmp894 = mem_1[tmp862];
    assign tmp620 = {tmp604, tmp609, tmp614, tmp619, tmp608, tmp613, tmp618, tmp607, tmp612, tmp617, tmp606, tmp611, tmp616, tmp605, tmp610, tmp615};
    assign tmp1168 = tmp1184;
    assign tmp241 = {shifted_w39[8], shifted_w39[9], shifted_w39[10], shifted_w39[11], shifted_w39[12], shifted_w39[13], shifted_w39[14], shifted_w39[15]};
    assign tmp1785 = {temp_21[48], temp_21[49], temp_21[50], temp_21[51], temp_21[52], temp_21[53], temp_21[54], temp_21[55]};
    assign tmp2914 = {temp_36[0], temp_36[1], temp_36[2], temp_36[3], temp_36[4], temp_36[5], temp_36[6], temp_36[7]};
    assign tmp1955 = tmp1951 ^ tmp1954;
    assign tmp1841 = {const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0, const1840_0};
    assign tmp1345 = tmp1341 ^ tmp1344;
    assign tmp1501 = {temp_18[112], temp_18[113], temp_18[114], temp_18[115], temp_18[116], temp_18[117], temp_18[118], temp_18[119]};
    assign tmp83 = tmp82 ^ tmp58;
    assign tmp2110 = tmp2225;
    assign tmp561 = {temp_4[72], temp_4[73], temp_4[74], temp_4[75], temp_4[76], temp_4[77], temp_4[78], temp_4[79]};
        assign tmp1042 = mem_3[tmp922];
    assign tmp1537 = {tmp1536, tmp1502};
    assign tmp2252 = tmp2250 ^ tmp2251;
        assign tmp2933 = mem_1[tmp2901];
    assign tmp1321 = tmp1317 ^ tmp1320;
        assign tmp149 = mem_2[const148_6];
    assign tmp1200 = {temp_13[40], temp_13[41], temp_13[42], temp_13[43], temp_13[44], temp_13[45], temp_13[46], temp_13[47]};
    assign tmp1065 = {tmp1064[0], tmp1064[1], tmp1064[2], tmp1064[3], tmp1064[4], tmp1064[5], tmp1064[6], tmp1064[7]};
    assign tmp2953 = {temp_37[80], temp_37[81], temp_37[82], temp_37[83], temp_37[84], temp_37[85], temp_37[86], temp_37[87]};
        assign tmp1533 = mem_4[tmp1501];
    assign tmp1340 = {tmp1339, tmp1217};
    assign tmp787 = tmp785 ^ tmp786;
    assign tmp2084 = {temp_25[0], temp_25[1], temp_25[2], temp_25[3], temp_25[4], temp_25[5], temp_25[6], temp_25[7]};
    assign tmp551 = {tmp550[0], tmp550[1], tmp550[2], tmp550[3], tmp550[4], tmp550[5], tmp550[6], tmp550[7]};
    assign tmp1815 = tmp1908;
    assign tmp1730 = {temp_20[96], temp_20[97], temp_20[98], temp_20[99], temp_20[100], temp_20[101], temp_20[102], temp_20[103]};
    assign tmp569 = {temp_4[8], temp_4[9], temp_4[10], temp_4[11], temp_4[12], temp_4[13], temp_4[14], temp_4[15]};
    assign tmp1995 = tmp1993 ^ tmp1994;
    assign tmp1963 = tmp1959 ^ tmp1962;
    assign tmp919 = {temp_10[80], temp_10[81], temp_10[82], temp_10[83], temp_10[84], temp_10[85], temp_10[86], temp_10[87]};
        assign tmp750 = mem_4[tmp630];
    assign tmp330 = {temp_2[104], temp_2[105], temp_2[106], temp_2[107], temp_2[108], temp_2[109], temp_2[110], temp_2[111]};
        assign tmp2447 = mem_3[tmp2382];
    assign tmp2960 = {temp_37[24], temp_37[25], temp_37[26], temp_37[27], temp_37[28], temp_37[29], temp_37[30], temp_37[31]};
    assign tmp1075 = {tmp1074, tmp923};
    assign tmp103 = {rc1_w15, rc2_w15, rc3_w15, rc4_w15};
    assign tmp1327 = {const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0, const1326_0};
    assign tmp2756 = {const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0, const2755_0};
        assign tmp591 = mem_1[tmp559];
    assign tmp1442 = {temp_16[56], temp_16[57], temp_16[58], temp_16[59], temp_16[60], temp_16[61], temp_16[62], temp_16[63]};
    assign tmp61 = {tmp58[8], tmp58[9], tmp58[10], tmp58[11], tmp58[12], tmp58[13], tmp58[14], tmp58[15]};
    assign tmp1846 = {tmp1845, tmp1793};
    assign tmp1728 = {temp_20[112], temp_20[113], temp_20[114], temp_20[115], temp_20[116], temp_20[117], temp_20[118], temp_20[119]};
    assign tmp1424 = {tmp1423, tmp1220};
    assign tmp134 = {tmp133[24], tmp133[25], tmp133[26], tmp133[27], tmp133[28], tmp133[29], tmp133[30], tmp133[31]};
    assign tmp1237 = tmp1418;
    assign tmp2386 = {temp_30[64], temp_30[65], temp_30[66], temp_30[67], temp_30[68], temp_30[69], temp_30[70], temp_30[71]};
    assign expanded_key = tmp259;

    always @( posedge clk )
    begin
    end
endmodule

module tb();
    reg clk;
    reg [127:0] aes_key;
    reg [127:0] aes_plaintext;
    wire [127:0] aes_ciphertext;

    toplevel block(.aes_key(aes_key), .aes_plaintext(aes_plaintext), .aes_ciphertext(aes_ciphertext), .clk(clk));

    always
        #0.5 clk = ~clk;

    initial begin
        $dumpfile ("waveform.vcd");
        $dumpvars;

        clk = 0;
        aes_key = 128'd0;
        aes_plaintext = 128'd0;

        #2
        $finish;
    end
endmodule
