--- Verilog for the Counter ---
module toplevel(aes_plaintext, aes_key, aes_ciphertext, clk);
    input[127:0] aes_ciphertext;
    input[127:0] aes_key;
    input clk;
    output[127:0] aes_plaintext;

    wire[255:0] tmp675;
    wire[255:0] tmp1993;
    wire[255:0] tmp1061;
    wire[7:0] tmp966;
    wire[7:0] tmp168;
    wire[7:0] tmp1421;
    wire[255:0] tmp1996;
    wire[7:0] tmp592;
    wire[255:0] tmp1376;
    wire[7:0] tmp1070;
    wire[255:0] tmp853;
    wire[7:0] tmp169;
    wire[7:0] tmp1000;
    wire[7:0] tmp955;
    wire[255:0] tmp1064;
    wire[7:0] tmp280;
    wire[255:0] tmp376;
    wire[7:0] tmp170;
    wire[127:0] tmp559;
    wire[255:0] tmp1065;
    wire[7:0] tmp2006;
    wire[255:0] tmp645;
    wire[255:0] tmp1999;
    wire[255:0] tmp1528;
    wire[7:0] c1_w27;
    wire[7:0] c2_w27;
    wire[255:0] tmp854;
    wire[7:0] c3_w27;
    wire[7:0] c4_w27;
    wire[7:0] tmp793;
    wire[255:0] tmp2311;
    wire[255:0] tmp1069;
    wire[7:0] tmp63;
    wire[7:0] tmp243;
    wire[255:0] tmp2003;
    wire[7:0] tmp956;
    wire[127:0] tmp172;
    wire[127:0] tmp1010;
    wire[255:0] tmp1074;
    wire[127:0] tmp281;
    wire[7:0] tmp1388;
    wire[255:0] tmp1381;
    wire[31:0] concat_w3;
    wire[127:0] tmp173;
    wire[7:0] a4_w27;
    wire[255:0] tmp1072;
    wire[255:0] tmp595;
    wire[255:0] tmp2320;
    wire[255:0] tmp855;
    wire[127:0] tmp174;
    wire[255:0] tmp2007;
    wire[255:0] tmp1113;
    wire[255:0] tmp1385;
    wire[255:0] tmp2306;
    wire[255:0] tmp2008;
    wire[31:0] tmp175;
    wire[255:0] tmp1322;
    wire[255:0] tmp2009;
    wire[7:0] tmp957;
    wire[255:0] tmp1077;
    wire[31:0] xor_w27;
    wire[255:0] tmp1066;
    wire[7:0] rc1_w27;
    wire[7:0] rc2_w27;
    wire[7:0] tmp2284;
    wire[7:0] rc3_w27;
    wire[7:0] rc4_w27;
    wire[255:0] tmp648;
    wire[255:0] tmp1082;
    wire[7:0] const178_0;
    wire[7:0] tmp64;
    wire[255:0] tmp2323;
    wire[7:0] tmp244;
    wire[127:0] tmp1465;
    wire[255:0] tmp1080;
    wire[7:0] const130_0;
    wire[7:0] tmp1424;
    wire[255:0] tmp1063;
    wire[255:0] tmp1081;
    wire[7:0] const179_0;
    wire[31:0] tmp32;
    wire[7:0] tmp1679;
    wire[7:0] tmp958;
    wire[7:0] tmp162;
    wire[7:0] tmp746;
    wire[7:0] tmp1681;
    wire[7:0] tmp1682;
    wire[7:0] tmp747;
    wire[7:0] tmp1684;
    wire[255:0] tmp1772;
    wire[7:0] tmp1685;
    wire[255:0] tmp649;
    wire[7:0] tmp748;
    wire[7:0] tmp1687;
    wire[7:0] tmp283;
    wire[7:0] tmp1688;
    wire[7:0] tmp749;
    wire[255:0] tmp860;
    wire[7:0] tmp1690;
    wire[255:0] tmp2330;
    wire[255:0] tmp1116;
    wire[7:0] tmp750;
    wire[7:0] tmp1693;
    wire[255:0] tmp1374;
    wire[127:0] tmp1710;
    wire[7:0] tmp751;
    wire[7:0] tmp864;
    wire[127:0] tmp493;
    wire[7:0] tmp752;
    wire[255:0] tmp659;
    wire[7:0] tmp1047;
    wire[7:0] tmp65;
    wire[127:0] tmp1695;
    wire[7:0] tmp753;
    wire[7:0] tmp245;
    wire[7:0] tmp1739;
    wire[7:0] tmp754;
    wire[127:0] tmp1696;
    wire[255:0] tmp1303;
    wire[7:0] tmp755;
    wire[7:0] tmp797;
    wire[7:0] tmp404;
    wire[7:0] tmp2336;
    wire[255:0] tmp599;
    wire[127:0] temp_5;
    wire[7:0] tmp757;
    wire[255:0] tmp1328;
    wire[7:0] tmp1776;
    wire[127:0] tmp1698;
    wire[7:0] tmp2338;
    wire[7:0] b1_w31;
    wire[7:0] tmp759;
    wire[255:0] tmp1532;
    wire[7:0] tmp760;
    wire[7:0] tmp761;
    wire[127:0] tmp562;
    wire[7:0] tmp762;
    wire[7:0] tmp763;
    wire[7:0] tmp764;
    wire[7:0] tmp765;
    wire[7:0] tmp285;
    wire[7:0] tmp766;
    wire[7:0] tmp767;
    wire[31:0] shifted_w23;
    wire[7:0] tmp768;
    wire[127:0] tmp1466;
    wire[7:0] tmp769;
    wire[31:0] shifted_w35;
    wire[7:0] tmp770;
    wire[7:0] tmp771;
    wire[31:0] shifted_w11;
    wire[7:0] tmp772;
    wire[7:0] tmp773;
    wire[31:0] tmp141;
    wire[127:0] tmp790;
    wire[127:0] tmp774;
    wire[127:0] tmp1018;
    wire[7:0] tmp961;
    wire[7:0] tmp2344;
    wire[7:0] tmp120;
    wire[127:0] tmp1702;
    wire[255:0] tmp1067;
    wire[7:0] tmp2345;
    wire[7:0] c2_w39;
    wire[127:0] tmp775;
    wire[7:0] tmp2346;
    wire[7:0] tmp286;
    wire[127:0] temp_6;
    wire[7:0] c2_w23;
    wire[255:0] tmp2015;
    wire[255:0] tmp668;
    wire[255:0] tmp427;
    wire[127:0] tmp776;
    wire[7:0] const180_0;
    wire[255:0] tmp1122;
    wire[127:0] tmp1704;
    wire[7:0] b2_w31;
    wire[255:0] tmp1394;
    wire[255:0] tmp1068;
    wire[31:0] concat_w27;
    wire[255:0] tmp2082;
    wire[31:0] tmp181;
    wire[255:0] tmp461;
    wire[31:0] xor_w15;
    wire[127:0] tmp1705;
    wire[255:0] tmp2209;
    wire[31:0] tmp182;
    wire[127:0] tmp778;
    wire[255:0] tmp2020;
    wire[255:0] tmp1400;
    wire[31:0] tmp183;
    wire[7:0] b1_w35;
    wire[255:0] tmp1397;
    wire[31:0] tmp184;
    wire[31:0] substituted_w27;
    wire[255:0] tmp465;
    wire[7:0] tmp1689;
    wire[31:0] tmp185;
    wire[7:0] b1_w23;
    wire[255:0] tmp466;
    wire[31:0] tmp186;
    wire[7:0] tmp800;
    wire[127:0] tmp780;
    wire[255:0] tmp467;
    wire[127:0] tmp171;
    wire[7:0] a2_w31;
    wire[7:0] a3_w31;
    wire[7:0] tmp1340;
    wire[7:0] b2_w23;
    wire[7:0] tmp1227;
    wire[7:0] a4_w31;
    wire[7:0] tmp187;
    wire[7:0] tmp963;
    wire[255:0] tmp1402;
    wire[255:0] tmp472;
    wire[7:0] b3_w11;
    wire[127:0] temp_7;
    wire[255:0] tmp2025;
    wire[255:0] tmp1403;
    wire[255:0] tmp395;
    wire[7:0] tmp188;
    wire[7:0] tmp527;
    wire[7:0] tmp497;
    wire[255:0] tmp2027;
    wire[7:0] b4_w11;
    wire[255:0] tmp2028;
    wire[7:0] tmp2086;
    wire[127:0] tmp783;
    wire[7:0] tmp1412;
    wire[7:0] c4_w15;
    wire[255:0] tmp2029;
    wire[7:0] tmp801;
    wire[127:0] new_4;
    wire[255:0] tmp473;
    wire[7:0] tmp610;
    wire[255:0] tmp1406;
    wire[255:0] tmp474;
    wire[127:0] tmp1479;
    wire[127:0] tmp1712;
    wire[255:0] tmp1407;
    wire[255:0] tmp475;
    wire[255:0] tmp660;
    wire[31:0] shifted_w31;
    wire[255:0] tmp603;
    wire[31:0] tmp191;
    wire[7:0] tmp340;
    wire[255:0] tmp1409;
    wire[255:0] tmp2032;
    wire[255:0] tmp1410;
    wire[31:0] tmp131;
    wire[255:0] tmp655;
    wire[255:0] tmp480;
    wire[31:0] tmp206;
    wire[7:0] tmp1714;
    wire[255:0] tmp2314;
    wire[255:0] tmp1411;
    wire[127:0] tmp148;
    wire[7:0] b4_w31;
    wire[7:0] tmp192;
    wire[255:0] tmp478;
    wire[127:0] tmp1431;
    wire[7:0] tmp1716;
    wire[255:0] tmp687;
    wire[255:0] tmp1384;
    wire[127:0] temp_8;
    wire[255:0] tmp479;
    wire[7:0] tmp193;
    wire[127:0] tmp788;
    wire[255:0] tmp1305;
    wire[255:0] tmp656;
    wire[7:0] tmp1206;
    wire[255:0] tmp638;
    wire[127:0] temp_18;
    wire[255:0] tmp1152;
    wire[7:0] tmp1078;
    wire[7:0] tmp1271;
    wire[255:0] tmp1083;
    wire[7:0] tmp484;
    wire[255:0] tmp1084;
    wire[7:0] tmp499;
    wire[255:0] tmp2005;
    wire[255:0] tmp1085;
    wire[7:0] tmp1944;
    wire[7:0] c1_w11;
    wire[255:0] tmp1123;
    wire[255:0] tmp2004;
    wire[255:0] tmp1090;
    wire[7:0] tmp1094;
    wire[255:0] tmp397;
    wire[255:0] tmp1087;
    wire[7:0] tmp2220;
    wire[7:0] tmp658;
    wire[255:0] tmp1088;
    wire[255:0] tmp1177;
    wire[127:0] tmp1250;
    wire[255:0] tmp1089;
    wire[255:0] tmp1124;
    wire[7:0] tmp163;
    wire[255:0] tmp1382;
    wire[255:0] tmp1091;
    wire[255:0] tmp843;
    wire[255:0] tmp1383;
    wire[255:0] tmp1092;
    wire[255:0] tmp1093;
    wire[255:0] tmp1539;
    wire[255:0] tmp477;
    wire[7:0] rc3_w15;
    wire[7:0] tmp1433;
    wire[255:0] tmp1098;
    wire[7:0] tmp1102;
    wire[255:0] tmp1095;
    wire[7:0] c2_w11;
    wire[255:0] tmp1125;
    wire[255:0] tmp1096;
    wire[255:0] tmp1073;
    wire[255:0] tmp1097;
    wire[255:0] tmp1843;
    wire[255:0] tmp1099;
    wire[7:0] tmp2324;
    wire[255:0] tmp1100;
    wire[7:0] tmp2109;
    wire[255:0] tmp662;
    wire[255:0] tmp1101;
    wire[255:0] tmp688;
    wire[255:0] tmp608;
    wire[127:0] temp_10;
    wire[255:0] tmp1822;
    wire[7:0] tmp666;
    wire[255:0] tmp1106;
    wire[7:0] tmp1110;
    wire[255:0] tmp1103;
    wire[7:0] tmp1718;
    wire[7:0] tmp194;
    wire[255:0] tmp1075;
    wire[7:0] tmp1719;
    wire[127:0] tmp1482;
    wire[7:0] tmp2046;
    wire[255:0] tmp2039;
    wire[7:0] tmp1279;
    wire[7:0] tmp195;
    wire[255:0] tmp661;
    wire[255:0] tmp2318;
    wire[255:0] tmp2040;
    wire[7:0] tmp1721;
    wire[7:0] c1_w31;
    wire[7:0] tmp1280;
    wire[7:0] c2_w31;
    wire[7:0] c3_w31;
    wire[255:0] tmp1076;
    wire[7:0] c4_w31;
    wire[31:0] substituted_w31;
    wire[127:0] tmp196;
    wire[255:0] tmp2044;
    wire[7:0] tmp1281;
    wire[7:0] tmp1724;
    wire[255:0] tmp2045;
    wire[127:0] tmp197;
    wire[7:0] tmp1053;
    wire[7:0] tmp1282;
    wire[7:0] tmp1726;
    wire[255:0] tmp1153;
    wire[255:0] tmp2319;
    wire[127:0] tmp198;
    wire[7:0] tmp1274;
    wire[7:0] tmp1727;
    wire[255:0] tmp2047;
    wire[7:0] tmp952;
    wire[7:0] const101_4;
    wire[7:0] tmp341;
    wire[7:0] tmp1728;
    wire[127:0] tmp199;
    wire[255:0] tmp1387;
    wire[7:0] tmp1546;
    wire[7:0] tmp1729;
    wire[7:0] c1_w23;
    wire[255:0] tmp1359;
    wire[7:0] tmp1730;
    wire[7:0] c4_w11;
    wire[7:0] tmp1731;
    wire[255:0] tmp2218;
    wire[31:0] tmp200;
    wire[7:0] tmp1733;
    wire[255:0] tmp1854;
    wire[7:0] tmp1734;
    wire[7:0] tmp808;
    wire[7:0] tmp1735;
    wire[7:0] tmp2112;
    wire[31:0] xor_w31;
    wire[7:0] rc1_w31;
    wire[7:0] rc2_w31;
    wire[255:0] tmp1127;
    wire[7:0] rc3_w31;
    wire[7:0] c3_w11;
    wire[7:0] rc4_w31;
    wire[7:0] const201_8;
    wire[7:0] const203_0;
    wire[127:0] tmp202;
    wire[7:0] tmp342;
    wire[7:0] tmp1744;
    wire[255:0] tmp1748;
    wire[7:0] tmp296;
    wire[7:0] tmp2062;
    wire[255:0] tmp1745;
    wire[7:0] c4_w23;
    wire[7:0] tmp530;
    wire[255:0] tmp2219;
    wire[7:0] const204_0;
    wire[255:0] tmp611;
    wire[7:0] b1_w11;
    wire[255:0] tmp2057;
    wire[7:0] tmp2113;
    wire[31:0] concat_w31;
    wire[7:0] tmp996;
    wire[7:0] tmp1430;
    wire[255:0] tmp1749;
    wire[255:0] tmp2012;
    wire[255:0] tmp481;
    wire[255:0] tmp1104;
    wire[31:0] substituted_w11;
    wire[255:0] tmp482;
    wire[255:0] tmp1852;
    wire[7:0] tmp1415;
    wire[255:0] tmp1105;
    wire[255:0] tmp1392;
    wire[255:0] tmp483;
    wire[7:0] tmp1416;
    wire[255:0] tmp870;
    wire[31:0] tmp208;
    wire[255:0] tmp1107;
    wire[31:0] tmp209;
    wire[31:0] tmp207;
    wire[255:0] tmp1108;
    wire[255:0] tmp1179;
    wire[127:0] input_wire_8;
    wire[7:0] tmp492;
    wire[7:0] tmp1485;
    wire[255:0] tmp485;
    wire[127:0] new_8;
    wire[7:0] tmp1419;
    wire[7:0] a2_w35;
    wire[127:0] tmp177;
    wire[7:0] a3_w35;
    wire[7:0] tmp1420;
    wire[127:0] tmp1470;
    wire[7:0] tmp212;
    wire[7:0] tmp1118;
    wire[255:0] tmp1111;
    wire[255:0] tmp489;
    wire[7:0] tmp213;
    wire[255:0] tmp405;
    wire[255:0] tmp490;
    wire[255:0] tmp1576;
    wire[7:0] tmp794;
    wire[255:0] tmp491;
    wire[255:0] tmp1550;
    wire[7:0] tmp214;
    wire[7:0] tmp795;
    wire[7:0] tmp2115;
    wire[255:0] tmp1115;
    wire[7:0] tmp1856;
    wire[7:0] tmp796;
    wire[7:0] tmp215;
    wire[255:0] tmp1390;
    wire[127:0] tmp494;
    wire[255:0] tmp1117;
    wire[7:0] tmp345;
    wire[255:0] tmp2315;
    wire[7:0] tmp1427;
    wire[31:0] tmp216;
    wire[255:0] tmp1857;
    wire[7:0] tmp495;
    wire[7:0] tmp799;
    wire[255:0] tmp406;
    wire[7:0] tmp1126;
    wire[7:0] tmp1436;
    wire[7:0] tmp496;
    wire[7:0] tmp508;
    wire[7:0] b2_w35;
    wire[7:0] b3_w35;
    wire[7:0] tmp302;
    wire[7:0] b4_w35;
    wire[7:0] tmp217;
    wire[7:0] tmp1487;
    wire[255:0] tmp429;
    wire[7:0] tmp498;
    wire[7:0] tmp802;
    wire[7:0] tmp303;
    wire[7:0] tmp218;
    wire[7:0] tmp803;
    wire[7:0] tmp1432;
    wire[7:0] tmp500;
    wire[7:0] tmp346;
    wire[7:0] tmp804;
    wire[7:0] tmp219;
    wire[127:0] tmp73;
    wire[7:0] tmp501;
    wire[127:0] tmp787;
    wire[7:0] tmp805;
    wire[7:0] tmp1954;
    wire[7:0] tmp1434;
    wire[7:0] tmp502;
    wire[7:0] tmp2353;
    wire[7:0] tmp1041;
    wire[255:0] tmp663;
    wire[7:0] tmp2347;
    wire[7:0] tmp503;
    wire[7:0] tmp1488;
    wire[7:0] tmp2348;
    wire[7:0] tmp504;
    wire[255:0] tmp2325;
    wire[7:0] tmp2349;
    wire[7:0] tmp505;
    wire[7:0] tmp2350;
    wire[7:0] tmp347;
    wire[7:0] tmp506;
    wire[7:0] tmp1680;
    wire[127:0] tmp2351;
    wire[7:0] tmp507;
    wire[255:0] tmp846;
    wire[255:0] tmp1386;
    wire[255:0] tmp947;
    wire[7:0] tmp2354;
    wire[7:0] tmp2352;
    wire[255:0] tmp1155;
    wire[127:0] tmp324;
    wire[7:0] tmp509;
    wire[7:0] tmp2118;
    wire[7:0] tmp510;
    wire[255:0] tmp2326;
    wire[7:0] tmp737;
    wire[255:0] tmp1540;
    wire[127:0] tmp511;
    wire[7:0] tmp348;
    wire[7:0] tmp1042;
    wire[7:0] tmp2356;
    wire[7:0] const176_7;
    wire[7:0] a3_w39;
    wire[7:0] tmp512;
    wire[7:0] tmp1683;
    wire[7:0] tmp2357;
    wire[255:0] tmp410;
    wire[255:0] tmp871;
    wire[7:0] tmp513;
    wire[7:0] tmp2355;
    wire[7:0] tmp2358;
    wire[7:0] tmp618;
    wire[7:0] tmp514;
    wire[7:0] tmp240;
    wire[7:0] tmp2359;
    wire[7:0] tmp2119;
    wire[7:0] tmp515;
    wire[7:0] tmp2360;
    wire[7:0] tmp516;
    wire[255:0] tmp2327;
    wire[7:0] tmp2361;
    wire[7:0] tmp517;
    wire[7:0] tmp349;
    wire[7:0] tmp2362;
    wire[7:0] tmp518;
    wire[7:0] tmp1686;
    wire[7:0] tmp2363;
    wire[255:0] tmp411;
    wire[7:0] tmp519;
    wire[7:0] tmp350;
    wire[7:0] tmp2364;
    wire[7:0] tmp520;
    wire[127:0] tmp222;
    wire[127:0] tmp1251;
    wire[7:0] tmp2365;
    wire[7:0] tmp1491;
    wire[7:0] tmp521;
    wire[7:0] tmp351;
    wire[7:0] tmp2366;
    wire[7:0] tmp522;
    wire[7:0] tmp2367;
    wire[7:0] tmp806;
    wire[7:0] tmp352;
    wire[255:0] tmp2060;
    wire[255:0] tmp1130;
    wire[255:0] tmp2329;
    wire[7:0] tmp1134;
    wire[255:0] tmp1751;
    wire[7:0] c1_w35;
    wire[7:0] c2_w35;
    wire[255:0] tmp1128;
    wire[7:0] c4_w35;
    wire[7:0] tmp809;
    wire[7:0] tmp1438;
    wire[7:0] tmp1492;
    wire[7:0] tmp1760;
    wire[255:0] tmp1753;
    wire[7:0] tmp1439;
    wire[255:0] tmp1131;
    wire[7:0] tmp1691;
    wire[255:0] tmp2064;
    wire[255:0] tmp1132;
    wire[7:0] tmp43;
    wire[127:0] tmp96;
    wire[255:0] tmp1750;
    wire[255:0] tmp2065;
    wire[7:0] tmp355;
    wire[255:0] tmp1133;
    wire[7:0] tmp820;
    wire[7:0] tmp1692;
    wire[7:0] tmp821;
    wire[7:0] tmp1442;
    wire[7:0] tmp1959;
    wire[7:0] tmp823;
    wire[255:0] tmp632;
    wire[255:0] tmp2068;
    wire[7:0] tmp356;
    wire[7:0] tmp1443;
    wire[7:0] tmp832;
    wire[255:0] tmp2010;
    wire[255:0] tmp1135;
    wire[7:0] tmp1444;
    wire[7:0] tmp1960;
    wire[7:0] rc4_w3;
    wire[255:0] tmp1136;
    wire[7:0] tmp1445;
    wire[255:0] tmp1129;
    wire[255:0] tmp2331;
    wire[255:0] tmp1181;
    wire[255:0] tmp1137;
    wire[255:0] tmp2056;
    wire[7:0] tmp1446;
    wire[7:0] tmp1961;
    wire[7:0] rc1_w35;
    wire[7:0] rc2_w35;
    wire[7:0] tmp358;
    wire[7:0] rc3_w35;
    wire[255:0] tmp1762;
    wire[127:0] tmp1694;
    wire[7:0] const226_9;
    wire[7:0] tmp1284;
    wire[7:0] tmp1448;
    wire[7:0] rc4_w23;
    wire[7:0] tmp1449;
    wire[255:0] tmp1141;
    wire[7:0] tmp359;
    wire[7:0] tmp1451;
    wire[7:0] tmp1452;
    wire[255:0] tmp1765;
    wire[7:0] tmp1454;
    wire[7:0] const151_6;
    wire[255:0] tmp1766;
    wire[7:0] const229_0;
    wire[7:0] tmp360;
    wire[7:0] tmp1150;
    wire[255:0] tmp833;
    wire[7:0] tmp1459;
    wire[7:0] tmp1460;
    wire[7:0] const153_0;
    wire[255:0] tmp1144;
    wire[127:0] tmp72;
    wire[7:0] tmp1462;
    wire[7:0] tmp361;
    wire[7:0] tmp1045;
    wire[7:0] tmp1463;
    wire[255:0] tmp835;
    wire[7:0] tmp2014;
    wire[255:0] tmp1769;
    wire[127:0] tmp152;
    wire[31:0] tmp232;
    wire[255:0] tmp1747;
    wire[255:0] tmp1147;
    wire[7:0] tmp362;
    wire[127:0] input_wire_7;
    wire[255:0] tmp2080;
    wire[255:0] tmp1148;
    wire[7:0] a4_w23;
    wire[7:0] tmp436;
    wire[255:0] tmp1771;
    wire[7:0] tmp363;
    wire[7:0] tmp165;
    wire[255:0] tmp640;
    wire[127:0] tmp2333;
    wire[255:0] tmp1773;
    wire[127:0] tmp1014;
    wire[255:0] tmp1774;
    wire[7:0] tmp364;
    wire[255:0] tmp1775;
    wire[127:0] tmp2334;
    wire[7:0] c4_w39;
    wire[127:0] tmp1700;
    wire[255:0] tmp1780;
    wire[7:0] tmp1784;
    wire[255:0] tmp1777;
    wire[7:0] a2_w7;
    wire[7:0] const255_0;
    wire[7:0] tmp372;
    wire[255:0] tmp1778;
    wire[255:0] tmp665;
    wire[255:0] tmp1779;
    wire[7:0] rc2_w23;
    wire[7:0] a3_w7;
    wire[255:0] tmp1590;
    wire[31:0] tmp135;
    wire[255:0] tmp1781;
    wire[255:0] tmp1782;
    wire[7:0] a4_w7;
    wire[127:0] tmp1473;
    wire[255:0] tmp1783;
    wire[7:0] tmp698;
    wire[7:0] tmp37;
    wire[255:0] tmp431;
    wire[255:0] tmp1788;
    wire[7:0] tmp1792;
    wire[255:0] tmp1785;
    wire[255:0] tmp1313;
    wire[255:0] tmp2239;
    wire[255:0] tmp1786;
    wire[7:0] const104_0;
    wire[255:0] tmp366;
    wire[7:0] tmp2335;
    wire[255:0] tmp1787;
    wire[255:0] tmp1329;
    wire[127:0] tmp1469;
    wire[255:0] tmp1789;
    wire[255:0] tmp1287;
    wire[255:0] tmp1790;
    wire[7:0] tmp299;
    wire[7:0] tmp815;
    wire[127:0] tmp247;
    wire[255:0] tmp1791;
    wire[255:0] tmp1588;
    wire[31:0] tmp210;
    wire[255:0] tmp1330;
    wire[7:0] tmp1800;
    wire[255:0] tmp367;
    wire[127:0] temp_36;
    wire[127:0] tmp1697;
    wire[127:0] temp_37;
    wire[127:0] temp_38;
    wire[255:0] tmp710;
    wire[127:0] temp_39;
    wire[255:0] tmp950;
    wire[1407:0] expanded_key;
    wire[31:0] tmp8;
    wire[31:0] tmp9;
    wire[31:0] tmp10;
    wire[31:0] tmp11;
    wire[7:0] a1_w3;
    wire[7:0] a1_w27;
    wire[7:0] a2_w3;
    wire[255:0] tmp2235;
    wire[7:0] a3_w3;
    wire[7:0] tmp2378;
    wire[7:0] tmp12;
    wire[7:0] tmp2380;
    wire[255:0] tmp1641;
    wire[7:0] tmp528;
    wire[7:0] tmp529;
    wire[7:0] tmp13;
    wire[7:0] tmp531;
    wire[7:0] tmp2337;
    wire[7:0] tmp532;
    wire[7:0] tmp300;
    wire[7:0] tmp533;
    wire[7:0] tmp816;
    wire[127:0] tmp248;
    wire[7:0] tmp534;
    wire[7:0] tmp1054;
    wire[7:0] tmp535;
    wire[7:0] tmp536;
    wire[7:0] tmp537;
    wire[7:0] tmp538;
    wire[7:0] tmp539;
    wire[255:0] tmp868;
    wire[7:0] tmp15;
    wire[7:0] tmp541;
    wire[7:0] tmp542;
    wire[7:0] tmp543;
    wire[127:0] tmp560;
    wire[127:0] tmp544;
    wire[7:0] tmp39;
    wire[31:0] tmp16;
    wire[127:0] tmp1472;
    wire[255:0] tmp370;
    wire[7:0] tmp758;
    wire[7:0] b1_w3;
    wire[7:0] b2_w3;
    wire[255:0] tmp1799;
    wire[127:0] tmp2388;
    wire[7:0] b4_w3;
    wire[7:0] tmp17;
    wire[127:0] tmp546;
    wire[255:0] tmp1543;
    wire[127:0] tmp1474;
    wire[7:0] tmp18;
    wire[255:0] tmp2240;
    wire[127:0] tmp547;
    wire[127:0] tmp1475;
    wire[7:0] tmp301;
    wire[255:0] tmp1336;
    wire[7:0] tmp19;
    wire[127:0] tmp548;
    wire[255:0] tmp371;
    wire[127:0] tmp1021;
    wire[127:0] tmp1476;
    wire[7:0] tmp2339;
    wire[7:0] tmp20;
    wire[7:0] tmp2094;
    wire[255:0] tmp1176;
    wire[127:0] tmp549;
    wire[127:0] tmp1477;
    wire[7:0] tmp1086;
    wire[127:0] tmp1699;
    wire[7:0] c1_w3;
    wire[127:0] tmp550;
    wire[7:0] rc3_w39;
    wire[31:0] tmp233;
    wire[255:0] tmp2081;
    wire[31:0] substituted_w3;
    wire[127:0] tmp21;
    wire[31:0] tmp235;
    wire[255:0] tmp2083;
    wire[31:0] tmp236;
    wire[7:0] tmp1901;
    wire[255:0] tmp2084;
    wire[255:0] tmp844;
    wire[7:0] tmp2340;
    wire[7:0] tmp1158;
    wire[255:0] tmp841;
    wire[255:0] tmp867;
    wire[7:0] a4_w39;
    wire[7:0] tmp237;
    wire[7:0] tmp1435;
    wire[127:0] tmp23;
    wire[127:0] tmp553;
    wire[255:0] tmp2090;
    wire[7:0] tmp818;
    wire[31:0] tmp250;
    wire[7:0] tmp238;
    wire[255:0] tmp2087;
    wire[127:0] tmp554;
    wire[255:0] tmp845;
    wire[255:0] tmp2088;
    wire[7:0] tmp137;
    wire[7:0] tmp239;
    wire[31:0] tmp25;
    wire[255:0] tmp2089;
    wire[7:0] tmp807;
    wire[255:0] tmp847;
    wire[255:0] tmp1079;
    wire[127:0] tmp2398;
    wire[7:0] tmp2341;
    wire[31:0] xor_w3;
    wire[7:0] rc1_w3;
    wire[127:0] tmp1019;
    wire[127:0] tmp556;
    wire[7:0] rc3_w3;
    wire[255:0] tmp2061;
    wire[255:0] tmp1162;
    wire[31:0] shifted_w39;
    wire[7:0] b3_w39;
    wire[7:0] const28_0;
    wire[127:0] tmp27;
    wire[31:0] tmp41;
    wire[255:0] tmp850;
    wire[7:0] b1_w39;
    wire[7:0] b2_w39;
    wire[255:0] tmp851;
    wire[7:0] b4_w39;
    wire[255:0] tmp1802;
    wire[7:0] const29_0;
    wire[127:0] new_1;
    wire[7:0] tmp1903;
    wire[255:0] tmp1163;
    wire[7:0] const30_0;
    wire[7:0] tmp2342;
    wire[255:0] tmp1164;
    wire[127:0] tmp2402;
    wire[7:0] tmp819;
    wire[7:0] rc1_w39;
    wire[255:0] tmp2097;
    wire[31:0] tmp31;
    wire[7:0] c3_w35;
    wire[255:0] tmp2099;
    wire[127:0] input_wire_9;
    wire[255:0] tmp2100;
    wire[255:0] tmp1170;
    wire[7:0] rc2_w15;
    wire[127:0] tmp557;
    wire[127:0] new_9;
    wire[31:0] tmp33;
    wire[127:0] tmp1701;
    wire[127:0] temp_25;
    wire[31:0] tmp34;
    wire[255:0] tmp1803;
    wire[7:0] tmp856;
    wire[255:0] tmp858;
    wire[7:0] tmp1396;
    wire[31:0] tmp35;
    wire[31:0] substituted_w35;
    wire[7:0] c1_w39;
    wire[255:0] tmp859;
    wire[7:0] tmp2343;
    wire[127:0] tmp2104;
    wire[7:0] rc4_w39;
    wire[127:0] tmp1478;
    wire[127:0] tmp221;
    wire[255:0] tmp951;
    wire[7:0] tmp307;
    wire[7:0] tmp2105;
    wire[7:0] const251_10;
    wire[7:0] tmp2070;
    wire[7:0] tmp2106;
    wire[7:0] tmp2107;
    wire[7:0] const253_0;
    wire[127:0] input_wire_5;
    wire[7:0] tmp812;
    wire[7:0] tmp2108;
    wire[127:0] new_5;
    wire[127:0] tmp1481;
    wire[127:0] tmp252;
    wire[7:0] tmp739;
    wire[7:0] tmp813;
    wire[7:0] tmp2110;
    wire[127:0] temp_26;
    wire[7:0] tmp2111;
    wire[255:0] tmp715;
    wire[255:0] tmp849;
    wire[255:0] tmp434;
    wire[255:0] tmp1389;
    wire[7:0] tmp814;
    wire[7:0] tmp1483;
    wire[7:0] tmp1484;
    wire[255:0] tmp1756;
    wire[255:0] tmp1754;
    wire[7:0] tmp2114;
    wire[7:0] tmp1048;
    wire[7:0] tmp1486;
    wire[255:0] tmp876;
    wire[7:0] tmp1440;
    wire[7:0] tmp2116;
    wire[7:0] tmp674;
    wire[7:0] tmp2117;
    wire[127:0] tmp1184;
    wire[7:0] b3_w15;
    wire[7:0] tmp817;
    wire[7:0] tmp1489;
    wire[7:0] tmp1490;
    wire[255:0] tmp596;
    wire[255:0] tmp1807;
    wire[255:0] tmp1755;
    wire[7:0] tmp2120;
    wire[127:0] tmp1703;
    wire[127:0] tmp2121;
    wire[255:0] tmp1621;
    wire[127:0] tmp1022;
    wire[7:0] tmp1441;
    wire[7:0] tmp1493;
    wire[7:0] tmp2122;
    wire[7:0] tmp1166;
    wire[7:0] tmp1494;
    wire[255:0] tmp717;
    wire[7:0] tmp2123;
    wire[127:0] tmp223;
    wire[7:0] c3_w39;
    wire[7:0] a1_w7;
    wire[127:0] tmp741;
    wire[31:0] substituted_w39;
    wire[255:0] tmp861;
    wire[255:0] tmp1794;
    wire[255:0] tmp670;
    wire[255:0] tmp862;
    wire[255:0] tmp667;
    wire[255:0] tmp1795;
    wire[255:0] tmp863;
    wire[255:0] tmp1341;
    wire[7:0] tmp38;
    wire[7:0] b4_w15;
    wire[7:0] tmp822;
    wire[255:0] tmp1797;
    wire[7:0] a4_w35;
    wire[255:0] tmp1798;
    wire[255:0] tmp1178;
    wire[7:0] tmp44;
    wire[7:0] tmp1182;
    wire[255:0] tmp2066;
    wire[255:0] tmp1175;
    wire[255:0] tmp486;
    wire[7:0] const105_0;
    wire[127:0] tmp249;
    wire[255:0] tmp1393;
    wire[255:0] tmp866;
    wire[127:0] temp_28;
    wire[7:0] tmp40;
    wire[255:0] tmp1812;
    wire[255:0] tmp1804;
    wire[255:0] tmp1758;
    wire[7:0] tmp1808;
    wire[255:0] tmp1801;
    wire[255:0] tmp2016;
    wire[255:0] tmp1159;
    wire[31:0] shifted_w7;
    wire[255:0] tmp869;
    wire[255:0] tmp1342;
    wire[31:0] xor_w39;
    wire[255:0] tmp1180;
    wire[127:0] tmp224;
    wire[7:0] rc2_w39;
    wire[7:0] b1_w7;
    wire[7:0] tmp309;
    wire[7:0] b2_w7;
    wire[255:0] tmp415;
    wire[7:0] b3_w7;
    wire[31:0] concat_w39;
    wire[7:0] b4_w7;
    wire[7:0] tmp42;
    wire[7:0] tmp1913;
    wire[255:0] tmp1058;
    wire[255:0] tmp1806;
    wire[255:0] tmp464;
    wire[127:0] tmp1183;
    wire[7:0] tmp880;
    wire[255:0] tmp873;
    wire[255:0] tmp825;
    wire[7:0] const254_0;
    wire[255:0] tmp874;
    wire[7:0] tmp468;
    wire[7:0] tmp1185;
    wire[7:0] tmp1032;
    wire[7:0] tmp45;
    wire[255:0] tmp875;
    wire[7:0] tmp1816;
    wire[7:0] tmp1186;
    wire[31:0] tmp256;
    wire[7:0] tmp650;
    wire[255:0] tmp1395;
    wire[255:0] tmp877;
    wire[127:0] temp_29;
    wire[7:0] tmp1187;
    wire[127:0] tmp791;
    wire[255:0] tmp1810;
    wire[255:0] tmp878;
    wire[255:0] tmp435;
    wire[31:0] tmp257;
    wire[7:0] tmp1916;
    wire[7:0] tmp1188;
    wire[255:0] tmp879;
    wire[7:0] tmp313;
    wire[7:0] c2_w7;
    wire[31:0] tmp258;
    wire[255:0] tmp1813;
    wire[31:0] tmp259;
    wire[31:0] tmp225;
    wire[255:0] tmp1805;
    wire[127:0] tmp46;
    wire[31:0] tmp260;
    wire[127:0] tmp330;
    wire[7:0] tmp888;
    wire[7:0] tmp1208;
    wire[31:0] tmp261;
    wire[7:0] tmp1025;
    wire[7:0] tmp1918;
    wire[127:0] tmp47;
    wire[255:0] tmp1855;
    wire[7:0] tmp563;
    wire[255:0] tmp462;
    wire[255:0] tmp2011;
    wire[7:0] tmp2125;
    wire[255:0] tmp1811;
    wire[255:0] tmp1820;
    wire[7:0] tmp1824;
    wire[255:0] tmp1817;
    wire[7:0] tmp565;
    wire[7:0] tmp242;
    wire[255:0] tmp1818;
    wire[7:0] c1_w7;
    wire[127:0] tmp49;
    wire[255:0] tmp827;
    wire[255:0] tmp1819;
    wire[7:0] b2_w27;
    wire[7:0] tmp567;
    wire[255:0] tmp643;
    wire[127:0] temp_30;
    wire[31:0] tmp50;
    wire[7:0] tmp1655;
    wire[255:0] tmp1821;
    wire[7:0] tmp1717;
    wire[127:0] tmp953;
    wire[31:0] xor_w35;
    wire[7:0] tmp2130;
    wire[31:0] xor_w7;
    wire[255:0] tmp463;
    wire[7:0] rc1_w7;
    wire[7:0] tmp2131;
    wire[7:0] c3_w7;
    wire[255:0] tmp382;
    wire[7:0] rc3_w7;
    wire[7:0] rc4_w7;
    wire[255:0] tmp1761;
    wire[7:0] const51_2;
    wire[7:0] tmp571;
    wire[7:0] tmp1404;
    wire[127:0] tmp52;
    wire[255:0] tmp1607;
    wire[255:0] tmp1828;
    wire[7:0] c4_w7;
    wire[7:0] tmp572;
    wire[255:0] tmp1825;
    wire[7:0] tmp1923;
    wire[7:0] tmp2134;
    wire[255:0] tmp1055;
    wire[7:0] tmp573;
    wire[255:0] tmp2021;
    wire[255:0] tmp1826;
    wire[7:0] const54_0;
    wire[7:0] tmp140;
    wire[31:0] substituted_w7;
    wire[7:0] tmp574;
    wire[255:0] tmp1827;
    wire[255:0] tmp829;
    wire[7:0] const55_0;
    wire[7:0] tmp575;
    wire[127:0] tmp779;
    wire[31:0] concat_w7;
    wire[7:0] tmp1190;
    wire[7:0] tmp576;
    wire[255:0] tmp1830;
    wire[255:0] tmp487;
    wire[255:0] tmp2072;
    wire[7:0] tmp2138;
    wire[7:0] tmp577;
    wire[255:0] tmp1558;
    wire[31:0] tmp57;
    wire[7:0] tmp2141;
    wire[255:0] tmp884;
    wire[7:0] tmp578;
    wire[7:0] tmp2143;
    wire[255:0] tmp830;
    wire[7:0] c3_w19;
    wire[31:0] tmp58;
    wire[7:0] tmp579;
    wire[255:0] tmp1398;
    wire[255:0] tmp1160;
    wire[7:0] tmp580;
    wire[7:0] tmp581;
    wire[7:0] tmp1028;
    wire[31:0] tmp60;
    wire[7:0] tmp583;
    wire[7:0] const228_0;
    wire[31:0] tmp107;
    wire[31:0] tmp61;
    wire[7:0] tmp585;
    wire[7:0] a1_w11;
    wire[7:0] tmp587;
    wire[255:0] tmp881;
    wire[7:0] tmp588;
    wire[7:0] tmp589;
    wire[127:0] tmp227;
    wire[7:0] tmp590;
    wire[7:0] tmp591;
    wire[127:0] tmp316;
    wire[7:0] tmp1495;
    wire[7:0] rc2_w3;
    wire[1407:0] tmp262;
    wire[255:0] tmp882;
    wire[255:0] tmp831;
    wire[7:0] tmp1496;
    wire[255:0] tmp2321;
    wire[7:0] tmp810;
    wire[255:0] tmp1399;
    wire[127:0] new_state;
    wire[127:0] input_wire_11;
    wire[7:0] tmp725;
    wire[7:0] tmp1194;
    wire[127:0] tmp1925;
    wire[127:0] new_11;
    wire[127:0] tmp263;
    wire[7:0] a1_w31;
    wire[255:0] tmp886;
    wire[31:0] tmp133;
    wire[127:0] temp_32;
    wire[7:0] tmp848;
    wire[7:0] tmp1499;
    wire[7:0] tmp2124;
    wire[127:0] tmp264;
    wire[255:0] tmp1391;
    wire[7:0] tmp1501;
    wire[255:0] tmp678;
    wire[127:0] tmp1009;
    wire[7:0] tmp1502;
    wire[7:0] tmp1503;
    wire[127:0] tmp1708;
    wire[7:0] tmp1197;
    wire[7:0] tmp1505;
    wire[7:0] tmp265;
    wire[255:0] tmp892;
    wire[7:0] tmp1453;
    wire[7:0] tmp896;
    wire[7:0] tmp266;
    wire[7:0] tmp1199;
    wire[7:0] tmp1511;
    wire[7:0] tmp726;
    wire[255:0] tmp890;
    wire[7:0] tmp1200;
    wire[7:0] tmp1905;
    wire[7:0] tmp1514;
    wire[255:0] tmp891;
    wire[255:0] tmp1401;
    wire[7:0] tmp1522;
    wire[127:0] tmp777;
    wire[255:0] tmp1515;
    wire[7:0] tmp1030;
    wire[7:0] tmp269;
    wire[255:0] tmp893;
    wire[7:0] tmp1455;
    wire[7:0] tmp1202;
    wire[255:0] tmp894;
    wire[127:0] tmp781;
    wire[7:0] tmp1203;
    wire[7:0] tmp564;
    wire[255:0] tmp895;
    wire[255:0] tmp836;
    wire[7:0] tmp1204;
    wire[7:0] tmp167;
    wire[7:0] tmp272;
    wire[255:0] tmp644;
    wire[127:0] temp_33;
    wire[7:0] tmp1205;
    wire[127:0] tmp48;
    wire[7:0] tmp273;
    wire[7:0] a3_w11;
    wire[7:0] tmp904;
    wire[7:0] tmp840;
    wire[255:0] tmp1521;
    wire[7:0] tmp274;
    wire[127:0] tmp1709;
    wire[255:0] tmp898;
    wire[255:0] tmp1599;
    wire[7:0] tmp1031;
    wire[7:0] tmp275;
    wire[255:0] tmp1143;
    wire[255:0] tmp899;
    wire[7:0] tmp276;
    wire[7:0] tmp476;
    wire[255:0] tmp1523;
    wire[7:0] tmp1209;
    wire[255:0] tmp901;
    wire[255:0] tmp1524;
    wire[7:0] const230_0;
    wire[255:0] tmp902;
    wire[7:0] a1_w19;
    wire[7:0] tmp278;
    wire[255:0] tmp469;
    wire[255:0] tmp1525;
    wire[255:0] tmp903;
    wire[7:0] tmp728;
    wire[7:0] tmp279;
    wire[255:0] tmp677;
    wire[255:0] tmp2322;
    wire[127:0] tmp782;
    wire[127:0] tmp2155;
    wire[7:0] tmp2127;
    wire[255:0] tmp834;
    wire[127:0] tmp2156;
    wire[7:0] tmp566;
    wire[7:0] rc4_w11;
    wire[31:0] concat_w35;
    wire[127:0] tmp2157;
    wire[255:0] tmp470;
    wire[7:0] tmp729;
    wire[31:0] tmp231;
    wire[127:0] tmp2158;
    wire[7:0] tmp1554;
    wire[7:0] tmp2128;
    wire[255:0] tmp1367;
    wire[127:0] tmp2159;
    wire[255:0] tmp1145;
    wire[255:0] tmp2013;
    wire[127:0] tmp2160;
    wire[127:0] tmp1464;
    wire[7:0] tmp1024;
    wire[127:0] input_wire_4;
    wire[127:0] tmp2161;
    wire[255:0] tmp2079;
    wire[127:0] tmp558;
    wire[7:0] tmp1672;
    wire[127:0] tmp2162;
    wire[7:0] tmp2129;
    wire[255:0] tmp2226;
    wire[255:0] tmp2001;
    wire[127:0] tmp2163;
    wire[255:0] tmp1114;
    wire[255:0] tmp1405;
    wire[7:0] tmp568;
    wire[255:0] tmp837;
    wire[127:0] tmp2164;
    wire[7:0] tmp731;
    wire[127:0] tmp2165;
    wire[255:0] tmp1770;
    wire[255:0] tmp1860;
    wire[255:0] tmp1566;
    wire[255:0] tmp826;
    wire[127:0] tmp2166;
    wire[255:0] tmp838;
    wire[7:0] tmp190;
    wire[127:0] tmp2167;
    wire[7:0] tmp569;
    wire[255:0] tmp1815;
    wire[7:0] tmp1212;
    wire[7:0] tmp593;
    wire[7:0] tmp594;
    wire[255:0] tmp1563;
    wire[255:0] tmp598;
    wire[7:0] tmp602;
    wire[255:0] tmp1291;
    wire[255:0] tmp1529;
    wire[7:0] tmp1214;
    wire[7:0] tmp282;
    wire[7:0] tmp1215;
    wire[255:0] tmp1823;
    wire[255:0] tmp597;
    wire[7:0] tmp1216;
    wire[255:0] tmp1531;
    wire[7:0] tmp284;
    wire[255:0] tmp2034;
    wire[7:0] tmp1217;
    wire[255:0] tmp1842;
    wire[7:0] tmp570;
    wire[255:0] tmp600;
    wire[7:0] tmp1218;
    wire[31:0] tmp66;
    wire[255:0] tmp1057;
    wire[255:0] tmp601;
    wire[7:0] tmp2038;
    wire[7:0] tmp1221;
    wire[7:0] tmp1222;
    wire[7:0] tmp287;
    wire[7:0] b2_w11;
    wire[255:0] tmp1846;
    wire[7:0] tmp811;
    wire[7:0] tmp288;
    wire[127:0] tmp785;
    wire[7:0] tmp67;
    wire[7:0] tmp1228;
    wire[7:0] tmp2132;
    wire[7:0] tmp289;
    wire[7:0] tmp1230;
    wire[31:0] shifted_w19;
    wire[7:0] tmp1231;
    wire[7:0] tmp1418;
    wire[7:0] tmp1232;
    wire[7:0] tmp1233;
    wire[255:0] tmp1542;
    wire[7:0] const53_0;
    wire[127:0] tmp1234;
    wire[255:0] tmp1849;
    wire[255:0] tmp622;
    wire[31:0] tmp116;
    wire[7:0] tmp69;
    wire[255:0] tmp607;
    wire[255:0] tmp1565;
    wire[255:0] tmp1850;
    wire[127:0] tmp1235;
    wire[7:0] tmp293;
    wire[7:0] tmp70;
    wire[31:0] tmp109;
    wire[255:0] tmp609;
    wire[7:0] tmp294;
    wire[7:0] tmp1713;
    wire[127:0] tmp1236;
    wire[7:0] tmp744;
    wire[255:0] tmp1853;
    wire[7:0] tmp2133;
    wire[7:0] tmp295;
    wire[255:0] tmp1544;
    wire[127:0] tmp971;
    wire[255:0] tmp614;
    wire[127:0] tmp1237;
    wire[255:0] tmp671;
    wire[255:0] tmp1545;
    wire[127:0] tmp71;
    wire[7:0] tmp1832;
    wire[7:0] tmp297;
    wire[255:0] tmp612;
    wire[127:0] tmp1238;
    wire[7:0] tmp139;
    wire[255:0] tmp1154;
    wire[7:0] tmp298;
    wire[127:0] tmp786;
    wire[255:0] tmp613;
    wire[7:0] tmp1864;
    wire[255:0] tmp1138;
    wire[127:0] temp_3;
    wire[255:0] tmp1547;
    wire[255:0] tmp2063;
    wire[127:0] tmp1239;
    wire[255:0] tmp374;
    wire[255:0] tmp615;
    wire[7:0] tmp304;
    wire[255:0] tmp2033;
    wire[127:0] tmp1471;
    wire[7:0] tmp1039;
    wire[255:0] tmp908;
    wire[7:0] tmp912;
    wire[7:0] b3_w31;
    wire[255:0] tmp905;
    wire[7:0] tmp1437;
    wire[7:0] tmp1040;
    wire[7:0] tmp2140;
    wire[255:0] tmp906;
    wire[255:0] tmp1757;
    wire[7:0] tmp972;
    wire[127:0] temp_17;
    wire[255:0] tmp1568;
    wire[255:0] tmp907;
    wire[255:0] tmp1548;
    wire[7:0] tmp1257;
    wire[7:0] tmp1990;
    wire[7:0] b4_w19;
    wire[255:0] tmp909;
    wire[255:0] tmp828;
    wire[7:0] tmp1715;
    wire[255:0] tmp910;
    wire[7:0] tmp2135;
    wire[255:0] tmp911;
    wire[255:0] tmp2035;
    wire[255:0] tmp430;
    wire[7:0] tmp1027;
    wire[255:0] tmp2093;
    wire[255:0] tmp916;
    wire[7:0] tmp973;
    wire[7:0] tmp920;
    wire[255:0] tmp913;
    wire[255:0] tmp1569;
    wire[127:0] tmp2399;
    wire[127:0] temp_9;
    wire[255:0] tmp914;
    wire[255:0] tmp1601;
    wire[255:0] tmp915;
    wire[255:0] tmp2036;
    wire[7:0] tmp2136;
    wire[255:0] tmp917;
    wire[255:0] tmp918;
    wire[127:0] tmp1413;
    wire[7:0] rc4_w35;
    wire[7:0] tmp1046;
    wire[255:0] tmp919;
    wire[7:0] rc1_w23;
    wire[127:0] tmp1414;
    wire[255:0] tmp672;
    wire[7:0] tmp738;
    wire[255:0] tmp924;
    wire[7:0] tmp928;
    wire[7:0] tmp118;
    wire[255:0] tmp921;
    wire[255:0] tmp2037;
    wire[255:0] tmp922;
    wire[127:0] temp_13;
    wire[255:0] tmp923;
    wire[255:0] tmp2031;
    wire[255:0] tmp641;
    wire[31:0] tmp56;
    wire[255:0] tmp925;
    wire[7:0] tmp975;
    wire[7:0] tmp305;
    wire[255:0] tmp1112;
    wire[7:0] tmp306;
    wire[255:0] tmp1549;
    wire[7:0] tmp428;
    wire[127:0] temp_15;
    wire[7:0] tmp308;
    wire[255:0] tmp1371;
    wire[127:0] tmp2168;
    wire[255:0] tmp379;
    wire[7:0] tmp310;
    wire[7:0] tmp2178;
    wire[7:0] tmp311;
    wire[255:0] tmp616;
    wire[7:0] tmp312;
    wire[7:0] tmp745;
    wire[255:0] tmp1552;
    wire[255:0] tmp2067;
    wire[127:0] temp_16;
    wire[127:0] tmp2169;
    wire[127:0] tmp314;
    wire[255:0] tmp931;
    wire[255:0] tmp1553;
    wire[255:0] tmp1858;
    wire[255:0] tmp2018;
    wire[7:0] rc1_w11;
    wire[7:0] tmp2139;
    wire[127:0] tmp315;
    wire[7:0] tmp119;
    wire[127:0] input_wire_2;
    wire[7:0] tmp1026;
    wire[7:0] tmp1562;
    wire[127:0] tmp1240;
    wire[255:0] tmp1555;
    wire[127:0] new_2;
    wire[255:0] tmp1831;
    wire[127:0] tmp2171;
    wire[255:0] tmp1556;
    wire[127:0] tmp2172;
    wire[255:0] tmp617;
    wire[127:0] tmp317;
    wire[127:0] temp_19;
    wire[255:0] tmp1559;
    wire[7:0] tmp2173;
    wire[255:0] tmp1560;
    wire[7:0] tmp1213;
    wire[7:0] tmp2142;
    wire[7:0] tmp2174;
    wire[255:0] tmp1561;
    wire[127:0] tmp319;
    wire[7:0] tmp2175;
    wire[7:0] tmp1062;
    wire[7:0] tmp2176;
    wire[127:0] tmp320;
    wire[255:0] tmp664;
    wire[7:0] tmp722;
    wire[7:0] tmp1570;
    wire[7:0] rc3_w23;
    wire[7:0] tmp2177;
    wire[7:0] tmp2022;
    wire[127:0] temp_22;
    wire[255:0] tmp1564;
    wire[7:0] tmp388;
    wire[7:0] tmp2179;
    wire[127:0] tmp322;
    wire[7:0] tmp2145;
    wire[7:0] tmp2180;
    wire[255:0] tmp1567;
    wire[255:0] tmp381;
    wire[7:0] tmp2181;
    wire[127:0] tmp323;
    wire[31:0] tmp59;
    wire[7:0] tmp2182;
    wire[255:0] tmp1836;
    wire[7:0] tmp2183;
    wire[31:0] tmp75;
    wire[255:0] tmp1551;
    wire[7:0] tmp742;
    wire[7:0] tmp2144;
    wire[7:0] tmp526;
    wire[255:0] tmp926;
    wire[7:0] tmp1422;
    wire[255:0] tmp1809;
    wire[255:0] tmp1859;
    wire[7:0] tmp626;
    wire[255:0] tmp927;
    wire[127:0] tmp74;
    wire[7:0] tmp582;
    wire[255:0] tmp1861;
    wire[255:0] tmp2249;
    wire[127:0] tmp1241;
    wire[255:0] tmp1060;
    wire[255:0] tmp1862;
    wire[255:0] tmp619;
    wire[255:0] tmp932;
    wire[7:0] tmp936;
    wire[7:0] tmp2149;
    wire[255:0] tmp1863;
    wire[127:0] tmp1242;
    wire[31:0] xor_w11;
    wire[255:0] tmp2328;
    wire[255:0] tmp620;
    wire[7:0] rc2_w11;
    wire[7:0] tmp1189;
    wire[7:0] rc3_w11;
    wire[7:0] tmp584;
    wire[255:0] tmp621;
    wire[7:0] const76_3;
    wire[7:0] tmp2189;
    wire[7:0] c2_w19;
    wire[7:0] const78_0;
    wire[127:0] tmp77;
    wire[255:0] tmp623;
    wire[127:0] tmp1244;
    wire[255:0] tmp1834;
    wire[255:0] tmp934;
    wire[7:0] tmp980;
    wire[255:0] tmp1867;
    wire[7:0] tmp1840;
    wire[255:0] tmp625;
    wire[255:0] tmp930;
    wire[7:0] const79_0;
    wire[255:0] tmp1165;
    wire[7:0] tmp586;
    wire[255:0] tmp1869;
    wire[7:0] tmp1653;
    wire[7:0] const80_0;
    wire[255:0] tmp1759;
    wire[255:0] tmp1870;
    wire[255:0] tmp630;
    wire[7:0] tmp634;
    wire[255:0] tmp627;
    wire[7:0] a2_w11;
    wire[31:0] substituted_w19;
    wire[255:0] tmp2263;
    wire[255:0] tmp938;
    wire[31:0] tmp82;
    wire[255:0] tmp629;
    wire[127:0] tmp2170;
    wire[127:0] tmp1874;
    wire[31:0] tmp83;
    wire[127:0] tmp121;
    wire[7:0] tmp2332;
    wire[255:0] tmp941;
    wire[127:0] tmp1243;
    wire[255:0] tmp942;
    wire[7:0] a4_w11;
    wire[127:0] tmp1249;
    wire[31:0] tmp86;
    wire[7:0] tmp2190;
    wire[255:0] tmp943;
    wire[7:0] a1_w15;
    wire[7:0] tmp1872;
    wire[7:0] a2_w15;
    wire[255:0] tmp699;
    wire[7:0] a3_w15;
    wire[7:0] tmp62;
    wire[255:0] tmp1537;
    wire[7:0] a4_w15;
    wire[7:0] tmp87;
    wire[127:0] input_wire_6;
    wire[255:0] tmp1833;
    wire[7:0] tmp1878;
    wire[255:0] tmp1865;
    wire[255:0] tmp635;
    wire[127:0] new_6;
    wire[7:0] tmp1879;
    wire[7:0] tmp2146;
    wire[255:0] tmp946;
    wire[255:0] tmp386;
    wire[127:0] tmp1252;
    wire[7:0] tmp1914;
    wire[127:0] tmp325;
    wire[255:0] tmp933;
    wire[7:0] tmp1253;
    wire[255:0] tmp1527;
    wire[127:0] tmp326;
    wire[7:0] tmp1254;
    wire[127:0] tmp122;
    wire[255:0] tmp1866;
    wire[255:0] tmp1139;
    wire[7:0] tmp1255;
    wire[127:0] tmp327;
    wire[7:0] tmp1658;
    wire[255:0] tmp2098;
    wire[7:0] tmp1256;
    wire[7:0] tmp1723;
    wire[255:0] tmp387;
    wire[255:0] tmp624;
    wire[127:0] tmp328;
    wire[7:0] tmp1192;
    wire[7:0] tmp1258;
    wire[7:0] const154_0;
    wire[127:0] tmp329;
    wire[7:0] tmp1259;
    wire[7:0] tmp1610;
    wire[7:0] tmp2147;
    wire[7:0] tmp1260;
    wire[7:0] tmp1423;
    wire[7:0] tmp1261;
    wire[255:0] tmp2017;
    wire[127:0] input_wire_10;
    wire[255:0] tmp2069;
    wire[7:0] tmp1262;
    wire[127:0] new_10;
    wire[127:0] tmp331;
    wire[255:0] tmp935;
    wire[7:0] tmp1263;
    wire[7:0] tmp1892;
    wire[7:0] tmp1193;
    wire[127:0] tmp332;
    wire[7:0] tmp1264;
    wire[127:0] tmp123;
    wire[7:0] tmp1893;
    wire[127:0] tmp1245;
    wire[7:0] tmp1265;
    wire[7:0] tmp1894;
    wire[7:0] tmp1497;
    wire[7:0] tmp333;
    wire[255:0] tmp1541;
    wire[7:0] tmp1266;
    wire[7:0] tmp1895;
    wire[7:0] tmp334;
    wire[255:0] tmp1518;
    wire[7:0] tmp1267;
    wire[7:0] tmp1896;
    wire[255:0] tmp418;
    wire[7:0] tmp335;
    wire[7:0] tmp1268;
    wire[255:0] tmp392;
    wire[7:0] tmp1897;
    wire[7:0] tmp336;
    wire[7:0] tmp1269;
    wire[7:0] tmp1270;
    wire[7:0] tmp337;
    wire[7:0] tmp2148;
    wire[7:0] tmp1272;
    wire[7:0] tmp396;
    wire[7:0] tmp1899;
    wire[7:0] tmp338;
    wire[7:0] tmp1275;
    wire[7:0] tmp1276;
    wire[255:0] tmp885;
    wire[7:0] tmp339;
    wire[7:0] tmp1278;
    wire[7:0] tmp2184;
    wire[7:0] tmp89;
    wire[255:0] tmp419;
    wire[7:0] tmp2185;
    wire[255:0] tmp949;
    wire[127:0] tmp124;
    wire[255:0] tmp1837;
    wire[7:0] tmp90;
    wire[255:0] tmp940;
    wire[255:0] tmp1140;
    wire[7:0] tmp1195;
    wire[7:0] tmp2187;
    wire[7:0] tmp1447;
    wire[31:0] shifted_w15;
    wire[127:0] tmp561;
    wire[7:0] tmp2188;
    wire[7:0] tmp944;
    wire[127:0] input_wire_1;
    wire[255:0] tmp646;
    wire[7:0] b1_w15;
    wire[255:0] tmp390;
    wire[7:0] tmp2191;
    wire[255:0] tmp2301;
    wire[7:0] tmp2192;
    wire[255:0] tmp937;
    wire[7:0] b1_w19;
    wire[7:0] tmp2193;
    wire[255:0] tmp1994;
    wire[7:0] tmp92;
    wire[7:0] tmp1500;
    wire[7:0] tmp2195;
    wire[7:0] tmp2196;
    wire[7:0] tmp2197;
    wire[7:0] tmp2198;
    wire[7:0] tmp93;
    wire[7:0] tmp2200;
    wire[255:0] tmp887;
    wire[255:0] tmp647;
    wire[7:0] tmp2202;
    wire[7:0] tmp2203;
    wire[7:0] tmp94;
    wire[255:0] tmp2208;
    wire[7:0] tmp2212;
    wire[255:0] tmp2205;
    wire[7:0] tmp959;
    wire[31:0] tmp125;
    wire[7:0] tmp95;
    wire[255:0] tmp1151;
    wire[255:0] tmp2206;
    wire[255:0] tmp628;
    wire[7:0] tmp960;
    wire[255:0] tmp654;
    wire[255:0] tmp424;
    wire[255:0] tmp2207;
    wire[255:0] tmp651;
    wire[7:0] c2_w15;
    wire[7:0] c3_w15;
    wire[255:0] tmp652;
    wire[31:0] substituted_w15;
    wire[7:0] tmp1663;
    wire[255:0] tmp2210;
    wire[255:0] tmp653;
    wire[7:0] tmp989;
    wire[255:0] tmp2211;
    wire[7:0] tmp964;
    wire[127:0] tmp97;
    wire[255:0] tmp421;
    wire[255:0] tmp1323;
    wire[7:0] tmp2150;
    wire[7:0] tmp965;
    wire[255:0] tmp2216;
    wire[255:0] tmp939;
    wire[127:0] tmp98;
    wire[255:0] tmp2213;
    wire[7:0] tmp1498;
    wire[7:0] tmp1506;
    wire[255:0] tmp694;
    wire[7:0] tmp967;
    wire[255:0] tmp393;
    wire[255:0] tmp2214;
    wire[127:0] tmp99;
    wire[7:0] tmp968;
    wire[255:0] tmp2215;
    wire[7:0] tmp1198;
    wire[31:0] tmp36;
    wire[255:0] tmp1574;
    wire[7:0] tmp1578;
    wire[255:0] tmp1838;
    wire[255:0] tmp1571;
    wire[127:0] tmp1248;
    wire[255:0] tmp2217;
    wire[7:0] tmp1191;
    wire[7:0] tmp1283;
    wire[31:0] tmp158;
    wire[255:0] tmp1572;
    wire[255:0] tmp1288;
    wire[7:0] tmp523;
    wire[7:0] tmp1292;
    wire[255:0] tmp1573;
    wire[7:0] tmp343;
    wire[7:0] tmp1509;
    wire[255:0] tmp1286;
    wire[255:0] tmp857;
    wire[255:0] tmp1575;
    wire[7:0] tmp344;
    wire[255:0] tmp2224;
    wire[31:0] tmp84;
    wire[7:0] tmp2228;
    wire[255:0] tmp1357;
    wire[255:0] tmp2221;
    wire[7:0] tmp1665;
    wire[255:0] tmp1604;
    wire[255:0] tmp1577;
    wire[7:0] tmp2151;
    wire[255:0] tmp1289;
    wire[7:0] tmp2368;
    wire[255:0] tmp1764;
    wire[255:0] tmp2222;
    wire[255:0] tmp1290;
    wire[255:0] tmp2223;
    wire[255:0] tmp423;
    wire[255:0] tmp1582;
    wire[255:0] tmp883;
    wire[7:0] tmp1586;
    wire[7:0] tmp2369;
    wire[255:0] tmp1579;
    wire[255:0] tmp2225;
    wire[31:0] tmp85;
    wire[7:0] tmp682;
    wire[255:0] tmp1580;
    wire[7:0] tmp1512;
    wire[255:0] tmp1296;
    wire[7:0] tmp1300;
    wire[7:0] tmp2370;
    wire[255:0] tmp1293;
    wire[7:0] tmp353;
    wire[7:0] tmp1875;
    wire[7:0] tmp354;
    wire[255:0] tmp1294;
    wire[7:0] tmp1666;
    wire[255:0] tmp1583;
    wire[7:0] tmp357;
    wire[7:0] tmp2371;
    wire[255:0] tmp1295;
    wire[255:0] tmp2303;
    wire[7:0] tmp2236;
    wire[255:0] tmp2229;
    wire[255:0] tmp701;
    wire[255:0] tmp1585;
    wire[255:0] tmp1297;
    wire[255:0] tmp2230;
    wire[7:0] tmp2372;
    wire[31:0] concat_w11;
    wire[255:0] tmp1298;
    wire[255:0] tmp1835;
    wire[255:0] tmp368;
    wire[255:0] tmp633;
    wire[255:0] tmp2231;
    wire[7:0] tmp1174;
    wire[255:0] tmp1299;
    wire[7:0] tmp268;
    wire[7:0] tmp1594;
    wire[7:0] tmp2152;
    wire[255:0] tmp1587;
    wire[7:0] tmp2373;
    wire[7:0] tmp1768;
    wire[255:0] tmp2233;
    wire[7:0] tmp1876;
    wire[7:0] tmp1920;
    wire[255:0] tmp2234;
    wire[255:0] tmp1304;
    wire[127:0] tmp1201;
    wire[255:0] tmp1581;
    wire[7:0] tmp1308;
    wire[255:0] tmp1589;
    wire[7:0] tmp2374;
    wire[255:0] tmp369;
    wire[7:0] tmp1428;
    wire[255:0] tmp1302;
    wire[255:0] tmp1591;
    wire[255:0] tmp426;
    wire[255:0] tmp1349;
    wire[255:0] tmp1592;
    wire[127:0] tmp1467;
    wire[7:0] tmp2244;
    wire[7:0] tmp1029;
    wire[255:0] tmp2237;
    wire[255:0] tmp1593;
    wire[31:0] tmp100;
    wire[7:0] tmp2376;
    wire[7:0] tmp1902;
    wire[7:0] tmp1877;
    wire[7:0] tmp1429;
    wire[127:0] tmp2401;
    wire[255:0] tmp1598;
    wire[7:0] tmp1668;
    wire[7:0] rc1_w15;
    wire[255:0] tmp1595;
    wire[7:0] tmp2377;
    wire[31:0] tmp81;
    wire[7:0] tmp1904;
    wire[7:0] rc4_w15;
    wire[255:0] tmp1868;
    wire[255:0] tmp1596;
    wire[255:0] tmp1167;
    wire[7:0] const103_0;
    wire[255:0] tmp1516;
    wire[127:0] tmp102;
    wire[7:0] tmp2153;
    wire[255:0] tmp1597;
    wire[7:0] a4_w3;
    wire[7:0] tmp1425;
    wire[7:0] tmp1906;
    wire[255:0] tmp948;
    wire[7:0] tmp1907;
    wire[7:0] tmp270;
    wire[255:0] tmp2074;
    wire[255:0] tmp1763;
    wire[255:0] tmp1600;
    wire[7:0] tmp2379;
    wire[7:0] tmp1908;
    wire[7:0] tmp1909;
    wire[7:0] tmp642;
    wire[7:0] tmp1910;
    wire[127:0] tmp246;
    wire[7:0] tmp1911;
    wire[7:0] tmp1912;
    wire[31:0] concat_w15;
    wire[127:0] tmp1468;
    wire[31:0] tmp106;
    wire[255:0] tmp1839;
    wire[7:0] tmp1915;
    wire[255:0] tmp945;
    wire[255:0] tmp1606;
    wire[255:0] tmp1995;
    wire[7:0] tmp1917;
    wire[255:0] tmp1517;
    wire[255:0] tmp1603;
    wire[127:0] tmp1873;
    wire[7:0] tmp1919;
    wire[7:0] tmp2381;
    wire[7:0] tmp1450;
    wire[7:0] tmp1921;
    wire[31:0] tmp108;
    wire[7:0] tmp1196;
    wire[7:0] tmp271;
    wire[7:0] tmp2137;
    wire[255:0] tmp673;
    wire[7:0] tmp2382;
    wire[31:0] tmp110;
    wire[31:0] tmp156;
    wire[7:0] tmp88;
    wire[31:0] tmp111;
    wire[255:0] tmp1362;
    wire[255:0] tmp1605;
    wire[255:0] tmp1608;
    wire[7:0] tmp1656;
    wire[7:0] a2_w19;
    wire[7:0] tmp2383;
    wire[7:0] a3_w19;
    wire[7:0] a4_w19;
    wire[255:0] tmp636;
    wire[7:0] tmp1922;
    wire[7:0] tmp112;
    wire[127:0] tmp1926;
    wire[7:0] tmp2078;
    wire[255:0] tmp676;
    wire[127:0] tmp2400;
    wire[7:0] tmp1023;
    wire[7:0] tmp113;
    wire[127:0] tmp1927;
    wire[255:0] tmp1611;
    wire[255:0] tmp1519;
    wire[255:0] tmp365;
    wire[255:0] tmp679;
    wire[127:0] tmp2384;
    wire[255:0] tmp1612;
    wire[127:0] tmp1928;
    wire[7:0] tmp1880;
    wire[255:0] tmp1613;
    wire[255:0] tmp1363;
    wire[255:0] tmp681;
    wire[7:0] tmp115;
    wire[7:0] tmp2199;
    wire[7:0] tmp969;
    wire[255:0] tmp2238;
    wire[255:0] tmp1520;
    wire[7:0] tmp798;
    wire[7:0] tmp970;
    wire[7:0] tmp380;
    wire[255:0] tmp373;
    wire[255:0] tmp669;
    wire[255:0] tmp900;
    wire[255:0] tmp2241;
    wire[127:0] tmp2154;
    wire[127:0] tmp1020;
    wire[7:0] b2_w19;
    wire[7:0] tmp14;
    wire[255:0] tmp2242;
    wire[255:0] tmp375;
    wire[7:0] tmp117;
    wire[255:0] tmp2243;
    wire[127:0] tmp318;
    wire[255:0] tmp2071;
    wire[255:0] tmp377;
    wire[7:0] tmp974;
    wire[255:0] tmp378;
    wire[7:0] tmp1881;
    wire[7:0] tmp727;
    wire[255:0] tmp2248;
    wire[255:0] tmp897;
    wire[7:0] tmp2252;
    wire[7:0] tmp1380;
    wire[255:0] tmp2245;
    wire[127:0] tmp2385;
    wire[7:0] tmp976;
    wire[255:0] tmp2246;
    wire[7:0] tmp977;
    wire[255:0] tmp384;
    wire[255:0] tmp2247;
    wire[7:0] tmp978;
    wire[255:0] tmp2305;
    wire[255:0] tmp2042;
    wire[7:0] const155_0;
    wire[7:0] tmp979;
    wire[255:0] tmp1368;
    wire[7:0] c1_w19;
    wire[255:0] tmp2250;
    wire[255:0] tmp383;
    wire[7:0] c4_w19;
    wire[7:0] tmp1882;
    wire[255:0] tmp2251;
    wire[255:0] tmp1168;
    wire[7:0] tmp981;
    wire[7:0] tmp1207;
    wire[255:0] tmp385;
    wire[255:0] tmp2277;
    wire[7:0] tmp1142;
    wire[255:0] tmp1375;
    wire[7:0] tmp540;
    wire[7:0] tmp1426;
    wire[7:0] tmp982;
    wire[255:0] tmp1814;
    wire[127:0] tmp1940;
    wire[255:0] tmp2256;
    wire[7:0] tmp983;
    wire[255:0] tmp1365;
    wire[255:0] tmp2253;
    wire[7:0] tmp984;
    wire[255:0] tmp2254;
    wire[7:0] tmp1513;
    wire[7:0] tmp985;
    wire[255:0] tmp2255;
    wire[255:0] tmp389;
    wire[127:0] tmp2386;
    wire[255:0] tmp2227;
    wire[7:0] tmp986;
    wire[7:0] tmp1883;
    wire[255:0] tmp1847;
    wire[255:0] tmp2257;
    wire[7:0] tmp987;
    wire[255:0] tmp1526;
    wire[255:0] tmp2258;
    wire[255:0] tmp391;
    wire[7:0] tmp2201;
    wire[7:0] tmp988;
    wire[255:0] tmp2259;
    wire[7:0] tmp990;
    wire[7:0] tmp991;
    wire[7:0] tmp1530;
    wire[127:0] tmp1929;
    wire[7:0] tmp1223;
    wire[255:0] tmp1615;
    wire[255:0] tmp1616;
    wire[31:0] shifted_w27;
    wire[127:0] tmp1930;
    wire[255:0] tmp1617;
    wire[127:0] tmp1707;
    wire[31:0] shifted_w3;
    wire[7:0] tmp1884;
    wire[127:0] tmp1924;
    wire[255:0] tmp1609;
    wire[127:0] tmp1931;
    wire[255:0] tmp1622;
    wire[7:0] tmp1626;
    wire[255:0] tmp1619;
    wire[255:0] tmp2041;
    wire[127:0] tmp1932;
    wire[255:0] tmp1534;
    wire[7:0] tmp277;
    wire[255:0] tmp1620;
    wire[127:0] tmp2387;
    wire[127:0] tmp1933;
    wire[7:0] tmp1722;
    wire[255:0] tmp1146;
    wire[7:0] tmp1676;
    wire[7:0] c4_w3;
    wire[255:0] tmp1623;
    wire[255:0] tmp1630;
    wire[127:0] tmp1934;
    wire[255:0] tmp1624;
    wire[7:0] tmp1885;
    wire[7:0] tmp1210;
    wire[255:0] tmp1625;
    wire[127:0] tmp1935;
    wire[31:0] tmp157;
    wire[127:0] tmp1936;
    wire[7:0] tmp1634;
    wire[127:0] tmp545;
    wire[255:0] tmp1627;
    wire[255:0] tmp2043;
    wire[255:0] tmp1628;
    wire[255:0] tmp1369;
    wire[255:0] tmp1584;
    wire[255:0] tmp1629;
    wire[7:0] tmp1886;
    wire[127:0] tmp1938;
    wire[255:0] tmp1851;
    wire[7:0] tmp1538;
    wire[7:0] tmp1211;
    wire[255:0] tmp1631;
    wire[255:0] tmp1351;
    wire[7:0] b3_w3;
    wire[255:0] tmp1632;
    wire[127:0] tmp1939;
    wire[255:0] tmp1997;
    wire[7:0] b4_w27;
    wire[127:0] tmp1937;
    wire[255:0] tmp1638;
    wire[7:0] tmp444;
    wire[7:0] tmp1642;
    wire[255:0] tmp1635;
    wire[127:0] new_3;
    wire[127:0] tmp1941;
    wire[7:0] tmp1887;
    wire[7:0] b3_w19;
    wire[255:0] tmp1169;
    wire[7:0] rc1_w19;
    wire[7:0] tmp1219;
    wire[7:0] rc2_w19;
    wire[7:0] rc3_w19;
    wire[255:0] tmp2264;
    wire[7:0] tmp114;
    wire[7:0] tmp2268;
    wire[127:0] tmp1004;
    wire[255:0] tmp2261;
    wire[255:0] tmp1307;
    wire[7:0] tmp999;
    wire[255:0] tmp2262;
    wire[7:0] tmp1510;
    wire[7:0] tmp1001;
    wire[7:0] tmp1002;
    wire[7:0] tmp1725;
    wire[7:0] tmp1003;
    wire[255:0] tmp685;
    wire[127:0] tmp1246;
    wire[7:0] tmp1316;
    wire[255:0] tmp1309;
    wire[127:0] tmp2389;
    wire[255:0] tmp2265;
    wire[255:0] tmp1844;
    wire[7:0] tmp1888;
    wire[255:0] tmp2266;
    wire[127:0] tmp1005;
    wire[255:0] tmp929;
    wire[31:0] concat_w19;
    wire[255:0] tmp2267;
    wire[7:0] tmp2204;
    wire[255:0] tmp689;
    wire[7:0] tmp1456;
    wire[127:0] tmp1006;
    wire[255:0] tmp1171;
    wire[31:0] tmp132;
    wire[255:0] tmp1314;
    wire[7:0] tmp962;
    wire[31:0] xor_w19;
    wire[127:0] tmp1007;
    wire[255:0] tmp1315;
    wire[31:0] tmp134;
    wire[7:0] tmp1220;
    wire[255:0] tmp2270;
    wire[255:0] tmp692;
    wire[255:0] tmp1377;
    wire[127:0] tmp1008;
    wire[255:0] tmp2271;
    wire[7:0] tmp1889;
    wire[7:0] tmp189;
    wire[255:0] tmp693;
    wire[7:0] tmp1324;
    wire[7:0] a2_w23;
    wire[255:0] tmp2273;
    wire[255:0] tmp695;
    wire[255:0] tmp2274;
    wire[255:0] tmp2050;
    wire[255:0] tmp696;
    wire[255:0] tmp1319;
    wire[255:0] tmp1373;
    wire[255:0] tmp697;
    wire[127:0] tmp2390;
    wire[7:0] tmp138;
    wire[7:0] tmp1848;
    wire[7:0] tmp2054;
    wire[255:0] tmp1321;
    wire[127:0] tmp1011;
    wire[255:0] tmp1285;
    wire[255:0] tmp2280;
    wire[255:0] tmp702;
    wire[7:0] tmp706;
    wire[7:0] tmp1457;
    wire[255:0] tmp2307;
    wire[7:0] tmp1890;
    wire[127:0] tmp1012;
    wire[255:0] tmp2278;
    wire[255:0] tmp700;
    wire[255:0] tmp1327;
    wire[255:0] tmp2279;
    wire[127:0] tmp1013;
    wire[7:0] tmp1332;
    wire[255:0] tmp1325;
    wire[255:0] tmp2281;
    wire[255:0] tmp703;
    wire[255:0] tmp1633;
    wire[7:0] tmp2260;
    wire[255:0] tmp394;
    wire[127:0] tmp1942;
    wire[255:0] tmp2073;
    wire[7:0] b3_w23;
    wire[7:0] b4_w23;
    wire[31:0] tmp159;
    wire[7:0] tmp142;
    wire[127:0] tmp1891;
    wire[7:0] tmp1943;
    wire[255:0] tmp400;
    wire[127:0] tmp2391;
    wire[7:0] tmp143;
    wire[255:0] tmp1841;
    wire[7:0] tmp1945;
    wire[255:0] tmp398;
    wire[7:0] tmp2375;
    wire[7:0] tmp144;
    wire[7:0] tmp1946;
    wire[7:0] tmp1458;
    wire[255:0] tmp399;
    wire[255:0] tmp606;
    wire[255:0] tmp1172;
    wire[7:0] tmp1947;
    wire[7:0] tmp145;
    wire[255:0] tmp401;
    wire[7:0] tmp1948;
    wire[255:0] tmp402;
    wire[255:0] tmp2049;
    wire[255:0] tmp1119;
    wire[7:0] tmp1949;
    wire[255:0] tmp403;
    wire[7:0] c3_w23;
    wire[255:0] tmp1378;
    wire[7:0] tmp1950;
    wire[255:0] tmp2269;
    wire[31:0] substituted_w23;
    wire[127:0] tmp146;
    wire[7:0] tmp1951;
    wire[255:0] tmp2026;
    wire[255:0] tmp408;
    wire[7:0] tmp412;
    wire[127:0] input_wire_3;
    wire[255:0] tmp471;
    wire[7:0] tmp1952;
    wire[7:0] c1_w15;
    wire[127:0] tmp147;
    wire[7:0] tmp1732;
    wire[7:0] tmp1953;
    wire[127:0] tmp2392;
    wire[255:0] tmp2232;
    wire[255:0] tmp407;
    wire[7:0] tmp1955;
    wire[255:0] tmp409;
    wire[127:0] tmp149;
    wire[7:0] tmp1956;
    wire[255:0] tmp2051;
    wire[7:0] tmp1957;
    wire[31:0] tmp150;
    wire[7:0] tmp1958;
    wire[31:0] xor_w23;
    wire[255:0] tmp416;
    wire[255:0] tmp1557;
    wire[7:0] tmp420;
    wire[255:0] tmp413;
    wire[7:0] c2_w3;
    wire[7:0] tmp1962;
    wire[7:0] tmp1963;
    wire[255:0] tmp2052;
    wire[255:0] tmp414;
    wire[7:0] tmp1965;
    wire[7:0] tmp2030;
    wire[255:0] tmp1326;
    wire[255:0] tmp704;
    wire[7:0] tmp1737;
    wire[255:0] tmp1637;
    wire[7:0] tmp1964;
    wire[255:0] tmp705;
    wire[127:0] tmp1015;
    wire[7:0] c3_w3;
    wire[7:0] tmp68;
    wire[255:0] tmp1639;
    wire[7:0] tmp1738;
    wire[255:0] tmp1640;
    wire[127:0] tmp1016;
    wire[7:0] tmp756;
    wire[7:0] tmp714;
    wire[255:0] tmp2101;
    wire[255:0] tmp1331;
    wire[127:0] tmp2393;
    wire[127:0] tmp127;
    wire[255:0] tmp2053;
    wire[255:0] tmp708;
    wire[127:0] tmp1643;
    wire[31:0] tmp234;
    wire[127:0] tmp1644;
    wire[255:0] tmp1333;
    wire[7:0] tmp1740;
    wire[255:0] tmp711;
    wire[7:0] tmp1224;
    wire[255:0] tmp1334;
    wire[255:0] tmp712;
    wire[255:0] tmp422;
    wire[7:0] rc4_w19;
    wire[7:0] tmp1645;
    wire[7:0] tmp992;
    wire[255:0] tmp1335;
    wire[7:0] tmp1741;
    wire[255:0] tmp713;
    wire[7:0] tmp1646;
    wire[255:0] tmp2023;
    wire[255:0] tmp1636;
    wire[255:0] tmp1337;
    wire[7:0] const126_5;
    wire[7:0] tmp1647;
    wire[255:0] tmp1338;
    wire[7:0] tmp1742;
    wire[255:0] tmp718;
    wire[255:0] tmp680;
    wire[7:0] tmp1648;
    wire[127:0] tmp1247;
    wire[255:0] tmp1339;
    wire[127:0] new_7;
    wire[255:0] tmp2317;
    wire[7:0] const128_0;
    wire[7:0] tmp1649;
    wire[255:0] tmp716;
    wire[7:0] tmp1743;
    wire[7:0] tmp1650;
    wire[255:0] tmp2002;
    wire[255:0] tmp1344;
    wire[7:0] tmp1348;
    wire[127:0] tmp2394;
    wire[7:0] tmp1651;
    wire[7:0] tmp1461;
    wire[255:0] tmp719;
    wire[7:0] tmp1652;
    wire[255:0] tmp2048;
    wire[255:0] tmp720;
    wire[127:0] tmp22;
    wire[255:0] tmp1343;
    wire[127:0] tmp551;
    wire[255:0] tmp721;
    wire[255:0] tmp2058;
    wire[255:0] tmp1120;
    wire[7:0] tmp1654;
    wire[7:0] tmp1225;
    wire[255:0] tmp1345;
    wire[255:0] tmp839;
    wire[7:0] a1_w39;
    wire[255:0] tmp1346;
    wire[7:0] tmp993;
    wire[127:0] tmp723;
    wire[7:0] tmp1752;
    wire[127:0] tmp724;
    wire[255:0] tmp1347;
    wire[255:0] tmp2075;
    wire[127:0] tmp552;
    wire[7:0] tmp1657;
    wire[255:0] tmp1796;
    wire[255:0] tmp2055;
    wire[7:0] tmp1966;
    wire[255:0] tmp1533;
    wire[7:0] tmp1967;
    wire[7:0] tmp1968;
    wire[255:0] tmp2085;
    wire[7:0] tmp1969;
    wire[7:0] tmp1970;
    wire[7:0] tmp1971;
    wire[255:0] tmp707;
    wire[7:0] tmp290;
    wire[7:0] tmp1973;
    wire[7:0] tmp1974;
    wire[127:0] tmp2395;
    wire[255:0] tmp1978;
    wire[7:0] tmp1982;
    wire[7:0] tmp1898;
    wire[255:0] tmp1975;
    wire[255:0] tmp1173;
    wire[7:0] tmp1033;
    wire[255:0] tmp1976;
    wire[255:0] tmp1312;
    wire[7:0] tmp730;
    wire[7:0] tmp1034;
    wire[255:0] tmp1746;
    wire[255:0] tmp1977;
    wire[255:0] tmp1358;
    wire[255:0] tmp686;
    wire[7:0] tmp824;
    wire[7:0] tmp1226;
    wire[7:0] tmp1035;
    wire[7:0] rc2_w7;
    wire[255:0] tmp842;
    wire[255:0] tmp1979;
    wire[7:0] tmp994;
    wire[7:0] tmp1036;
    wire[255:0] tmp1980;
    wire[7:0] tmp733;
    wire[7:0] tmp1037;
    wire[255:0] tmp1981;
    wire[7:0] tmp734;
    wire[255:0] tmp1793;
    wire[127:0] temp_1;
    wire[7:0] tmp1273;
    wire[127:0] temp_2;
    wire[255:0] tmp2019;
    wire[7:0] tmp735;
    wire[127:0] temp_4;
    wire[255:0] tmp1986;
    wire[7:0] tmp736;
    wire[255:0] tmp1983;
    wire[7:0] const205_0;
    wire[7:0] tmp1043;
    wire[7:0] tmp1044;
    wire[255:0] tmp1984;
    wire[127:0] temp_11;
    wire[127:0] tmp2396;
    wire[127:0] temp_12;
    wire[255:0] tmp1985;
    wire[255:0] tmp2312;
    wire[255:0] tmp604;
    wire[127:0] temp_14;
    wire[7:0] tmp1050;
    wire[7:0] tmp1602;
    wire[7:0] tmp1051;
    wire[255:0] tmp1987;
    wire[255:0] tmp1310;
    wire[7:0] tmp740;
    wire[7:0] tmp1720;
    wire[255:0] tmp1988;
    wire[7:0] tmp1900;
    wire[127:0] temp_20;
    wire[7:0] tmp690;
    wire[127:0] temp_21;
    wire[7:0] tmp267;
    wire[255:0] tmp1989;
    wire[127:0] temp_23;
    wire[127:0] tmp24;
    wire[127:0] temp_24;
    wire[7:0] tmp995;
    wire[255:0] tmp1056;
    wire[7:0] tmp1277;
    wire[255:0] tmp631;
    wire[255:0] tmp1149;
    wire[127:0] temp_27;
    wire[255:0] tmp2024;
    wire[7:0] tmp743;
    wire[255:0] tmp2076;
    wire[255:0] tmp1379;
    wire[7:0] tmp1998;
    wire[255:0] tmp1991;
    wire[127:0] temp_31;
    wire[255:0] tmp2059;
    wire[255:0] tmp1059;
    wire[255:0] tmp1992;
    wire[127:0] temp_34;
    wire[127:0] temp_35;
    wire[255:0] tmp1311;
    wire[255:0] tmp2282;
    wire[7:0] tmp1504;
    wire[255:0] tmp1352;
    wire[7:0] tmp1356;
    wire[255:0] tmp2283;
    wire[255:0] tmp2313;
    wire[7:0] tmp1659;
    wire[127:0] tmp2397;
    wire[255:0] tmp417;
    wire[127:0] tmp1480;
    wire[255:0] tmp1350;
    wire[7:0] tmp2316;
    wire[255:0] tmp637;
    wire[7:0] tmp1660;
    wire[7:0] a2_w39;
    wire[255:0] tmp2288;
    wire[127:0] tmp1661;
    wire[255:0] tmp1156;
    wire[255:0] tmp2285;
    wire[31:0] concat_w23;
    wire[255:0] tmp1353;
    wire[255:0] tmp1121;
    wire[255:0] tmp683;
    wire[255:0] tmp2286;
    wire[255:0] tmp1354;
    wire[255:0] tmp1829;
    wire[7:0] tmp1049;
    wire[255:0] tmp2287;
    wire[255:0] tmp1767;
    wire[7:0] tmp524;
    wire[255:0] tmp1355;
    wire[7:0] tmp1972;
    wire[7:0] tmp1664;
    wire[255:0] tmp2289;
    wire[255:0] tmp889;
    wire[127:0] tmp555;
    wire[255:0] tmp2290;
    wire[255:0] tmp1360;
    wire[127:0] tmp789;
    wire[7:0] tmp1364;
    wire[255:0] tmp2291;
    wire[31:0] tmp161;
    wire[255:0] tmp425;
    wire[255:0] tmp1157;
    wire[7:0] tmp1667;
    wire[255:0] tmp1318;
    wire[7:0] a2_w27;
    wire[255:0] tmp639;
    wire[255:0] tmp2096;
    wire[7:0] a3_w27;
    wire[255:0] tmp2296;
    wire[7:0] tmp291;
    wire[7:0] tmp2300;
    wire[255:0] tmp2293;
    wire[255:0] tmp2272;
    wire[255:0] tmp1408;
    wire[7:0] tmp1669;
    wire[255:0] tmp1361;
    wire[255:0] tmp2309;
    wire[255:0] tmp2294;
    wire[7:0] tmp1670;
    wire[255:0] tmp432;
    wire[255:0] tmp1301;
    wire[255:0] tmp2295;
    wire[7:0] tmp2276;
    wire[7:0] tmp1671;
    wire[255:0] tmp2275;
    wire[7:0] tmp2186;
    wire[7:0] tmp164;
    wire[255:0] tmp2297;
    wire[7:0] tmp1229;
    wire[255:0] tmp1614;
    wire[31:0] tmp211;
    wire[255:0] tmp2298;
    wire[255:0] tmp2091;
    wire[7:0] tmp1673;
    wire[7:0] tmp997;
    wire[7:0] tmp1372;
    wire[255:0] tmp2299;
    wire[7:0] tmp1674;
    wire[255:0] tmp433;
    wire[255:0] tmp1306;
    wire[255:0] tmp1366;
    wire[127:0] tmp1711;
    wire[255:0] tmp691;
    wire[7:0] tmp1675;
    wire[31:0] tmp166;
    wire[255:0] tmp2304;
    wire[7:0] tmp2308;
    wire[255:0] tmp1535;
    wire[127:0] tmp784;
    wire[7:0] b1_w27;
    wire[255:0] tmp2092;
    wire[7:0] tmp1677;
    wire[7:0] b3_w27;
    wire[7:0] tmp1417;
    wire[255:0] tmp1370;
    wire[7:0] tmp1678;
    wire[255:0] tmp2000;
    wire[127:0] tmp2103;
    wire[255:0] tmp440;
    wire[7:0] tmp872;
    wire[255:0] tmp852;
    wire[255:0] tmp437;
    wire[255:0] tmp605;
    wire[255:0] tmp657;
    wire[255:0] tmp438;
    wire[7:0] tmp1662;
    wire[7:0] const26_1;
    wire[255:0] tmp439;
    wire[255:0] tmp488;
    wire[255:0] tmp1871;
    wire[255:0] tmp2302;
    wire[255:0] tmp441;
    wire[7:0] tmp1618;
    wire[31:0] tmp241;
    wire[255:0] tmp442;
    wire[7:0] tmp998;
    wire[7:0] tmp2292;
    wire[31:0] tmp91;
    wire[255:0] tmp443;
    wire[127:0] tmp321;
    wire[255:0] tmp2077;
    wire[7:0] tmp2126;
    wire[31:0] tmp136;
    wire[255:0] tmp1109;
    wire[255:0] tmp448;
    wire[7:0] tmp732;
    wire[7:0] tmp452;
    wire[255:0] tmp445;
    wire[255:0] tmp1320;
    wire[7:0] tmp1052;
    wire[7:0] tmp1507;
    wire[255:0] tmp446;
    wire[127:0] tmp1706;
    wire[255:0] tmp447;
    wire[255:0] tmp865;
    wire[7:0] a1_w23;
    wire[7:0] const129_0;
    wire[127:0] tmp1017;
    wire[7:0] a1_w35;
    wire[255:0] tmp449;
    wire[255:0] tmp450;
    wire[255:0] tmp1317;
    wire[127:0] tmp954;
    wire[255:0] tmp1071;
    wire[255:0] tmp451;
    wire[255:0] tmp684;
    wire[7:0] a3_w23;
    wire[7:0] tmp525;
    wire[7:0] b2_w15;
    wire[255:0] tmp456;
    wire[7:0] tmp460;
    wire[255:0] tmp453;
    wire[7:0] tmp1038;
    wire[255:0] tmp1161;
    wire[31:0] tmp160;
    wire[255:0] tmp454;
    wire[127:0] tmp792;
    wire[7:0] tmp220;
    wire[255:0] tmp1536;
    wire[255:0] tmp455;
    wire[7:0] tmp2102;
    wire[7:0] tmp1508;
    wire[255:0] tmp1845;
    wire[255:0] tmp457;
    wire[255:0] tmp709;
    wire[7:0] tmp292;
    wire[255:0] tmp458;
    wire[255:0] tmp2095;
    wire[7:0] tmp1736;
    wire[255:0] tmp459;
    wire[255:0] tmp2310;
    wire[7:0] tmp2194;

    reg[127:0] mem_2[255:0];
    reg[255:0] mem_6[255:0];
    reg[255:0] mem_7[255:0];
    reg[255:0] mem_5[255:0];
    reg[255:0] mem_4[255:0];
    reg[127:0] mem_1[255:0];
    reg[127:0] mem_3[255:0];

    assign const155_0 = 0;
    assign const251_10 = 10;
    assign const28_0 = 0;
    assign const180_0 = 0;
    assign const226_9 = 9;
    assign const126_5 = 5;
    assign const128_0 = 0;
    assign const55_0 = 0;
    assign const154_0 = 0;
    assign const26_1 = 1;
    assign const255_0 = 0;
    assign const228_0 = 0;
    assign const29_0 = 0;
    assign const101_4 = 4;
    assign const103_0 = 0;
    assign const253_0 = 0;
    assign const129_0 = 0;
    assign const201_8 = 8;
    assign const30_0 = 0;
    assign const203_0 = 0;
    assign const229_0 = 0;
    assign const105_0 = 0;
    assign const76_3 = 3;
    assign const54_0 = 0;
    assign const230_0 = 0;
    assign const104_0 = 0;
    assign const176_7 = 7;
    assign const178_0 = 0;
    assign const204_0 = 0;
    assign const78_0 = 0;
    assign const51_2 = 2;
    assign const53_0 = 0;
    assign const205_0 = 0;
    assign const130_0 = 0;
    assign const80_0 = 0;
    assign const79_0 = 0;
    assign const151_6 = 6;
    assign const254_0 = 0;
    assign const153_0 = 0;
    assign const179_0 = 0;
    assign tmp36 = tmp35 ^ tmp11;
        assign tmp1550 = mem_6[tmp1489];
    assign concat_w23 = tmp156;
        assign tmp1349 = mem_7[tmp1261];
    assign tmp387 = tmp385 ^ tmp386;
    assign tmp1134 = {tmp1133[0], tmp1133[1], tmp1133[2], tmp1133[3], tmp1133[4], tmp1133[5], tmp1133[6], tmp1133[7]};
    assign tmp232 = concat_w35 ^ substituted_w35;
    assign tmp1441 = {temp_21[48], temp_21[49], temp_21[50], temp_21[51], temp_21[52], temp_21[53], temp_21[54], temp_21[55]};
    assign rc3_w35 = const229_0;
        assign tmp1697 = mem_2[tmp1665];
    assign tmp540 = tmp556;
    assign tmp1259 = {temp_19[72], temp_19[73], temp_19[74], temp_19[75], temp_19[76], temp_19[77], temp_19[78], temp_19[79]};
    assign tmp1393 = tmp1391 ^ tmp1392;
        assign tmp2018 = mem_6[tmp1950];
        assign tmp1378 = mem_4[tmp1263];
    assign tmp1399 = tmp1397 ^ tmp1398;
    assign tmp1266 = {temp_19[16], temp_19[17], temp_19[18], temp_19[19], temp_19[20], temp_19[21], temp_19[22], temp_19[23]};
    assign tmp737 = {temp_8[24], temp_8[25], temp_8[26], temp_8[27], temp_8[28], temp_8[29], temp_8[30], temp_8[31]};
        assign tmp223 = mem_1[b3_w35];
    assign tmp344 = {temp_3[32], temp_3[33], temp_3[34], temp_3[35], temp_3[36], temp_3[37], temp_3[38], temp_3[39]};
    assign tmp615 = tmp613 ^ tmp614;
    assign tmp990 = tmp1006;
    assign tmp1674 = {temp_25[24], temp_25[25], temp_25[26], temp_25[27], temp_25[28], temp_25[29], temp_25[30], temp_25[31]};
    assign tmp363 = tmp484;
    assign tmp2361 = {temp_37[48], temp_37[49], temp_37[50], temp_37[51], temp_37[52], temp_37[53], temp_37[54], temp_37[55]};
        assign tmp1467 = mem_2[tmp1435];
    assign tmp1115 = tmp1113 ^ tmp1114;
    assign tmp1943 = {temp_31[120], temp_31[121], temp_31[122], temp_31[123], temp_31[124], temp_31[125], temp_31[126], temp_31[127]};
    assign tmp2127 = {temp_33[80], temp_33[81], temp_33[82], temp_33[83], temp_33[84], temp_33[85], temp_33[86], temp_33[87]};
    assign a1_w11 = tmp62;
    assign tmp1965 = tmp2030;
        assign tmp23 = mem_1[b3_w3];
    assign tmp1083 = tmp1081 ^ tmp1082;
    assign tmp1863 = tmp1861 ^ tmp1862;
        assign tmp1516 = mem_5[tmp1484];
    assign aes_plaintext = temp_39;
    assign tmp633 = tmp631 ^ tmp632;
        assign tmp643 = mem_7[tmp569];
        assign tmp1382 = mem_5[tmp1266];
        assign tmp1477 = mem_2[tmp1445];
    assign tmp1337 = tmp1335 ^ tmp1336;
        assign tmp2098 = mem_6[tmp1956];
    assign tmp2337 = {temp_36[104], temp_36[105], temp_36[106], temp_36[107], temp_36[108], temp_36[109], temp_36[110], temp_36[111]};
    assign tmp1890 = {temp_28[0], temp_28[1], temp_28[2], temp_28[3], temp_28[4], temp_28[5], temp_28[6], temp_28[7]};
    assign temp_25 = tmp1661;
    assign tmp1447 = {temp_21[0], temp_21[1], temp_21[2], temp_21[3], temp_21[4], temp_21[5], temp_21[6], temp_21[7]};
        assign tmp902 = mem_4[tmp801];
    assign tmp875 = tmp873 ^ tmp874;
        assign tmp247 = mem_1[b2_w39];
    assign tmp1279 = tmp1372;
        assign tmp1838 = mem_4[tmp1723];
    assign tmp1680 = tmp1696;
    assign concat_w39 = tmp256;
    assign a3_w31 = tmp189;
    assign tmp213 = {tmp211[16], tmp211[17], tmp211[18], tmp211[19], tmp211[20], tmp211[21], tmp211[22], tmp211[23]};
    assign temp_39 = new_1;
    assign tmp1982 = {tmp1981[0], tmp1981[1], tmp1981[2], tmp1981[3], tmp1981[4], tmp1981[5], tmp1981[6], tmp1981[7]};
    assign tmp2271 = tmp2269 ^ tmp2270;
    assign tmp275 = {new_state[40], new_state[41], new_state[42], new_state[43], new_state[44], new_state[45], new_state[46], new_state[47]};
        assign tmp554 = mem_2[tmp522];
    assign tmp168 = {shifted_w27[16], shifted_w27[17], shifted_w27[18], shifted_w27[19], shifted_w27[20], shifted_w27[21], shifted_w27[22], shifted_w27[23]};
    assign tmp2017 = tmp2015 ^ tmp2016;
    assign rc1_w3 = tmp27;
        assign tmp446 = mem_5[tmp344];
        assign tmp2039 = mem_7[tmp1951];
    assign tmp506 = {temp_4[32], temp_4[33], temp_4[34], temp_4[35], temp_4[36], temp_4[37], temp_4[38], temp_4[39]};
    assign tmp1881 = {temp_28[72], temp_28[73], temp_28[74], temp_28[75], temp_28[76], temp_28[77], temp_28[78], temp_28[79]};
        assign tmp624 = mem_4[tmp565];
    assign tmp108 = tmp83 ^ xor_w15;
    assign tmp579 = tmp602;
        assign tmp1828 = mem_6[tmp1721];
    assign tmp1711 = {expanded_key[896], expanded_key[897], expanded_key[898], expanded_key[899], expanded_key[900], expanded_key[901], expanded_key[902], expanded_key[903], expanded_key[904], expanded_key[905], expanded_key[906], expanded_key[907], expanded_key[908], expanded_key[909], expanded_key[910], expanded_key[911], expanded_key[912], expanded_key[913], expanded_key[914], expanded_key[915], expanded_key[916], expanded_key[917], expanded_key[918], expanded_key[919], expanded_key[920], expanded_key[921], expanded_key[922], expanded_key[923], expanded_key[924], expanded_key[925], expanded_key[926], expanded_key[927], expanded_key[928], expanded_key[929], expanded_key[930], expanded_key[931], expanded_key[932], expanded_key[933], expanded_key[934], expanded_key[935], expanded_key[936], expanded_key[937], expanded_key[938], expanded_key[939], expanded_key[940], expanded_key[941], expanded_key[942], expanded_key[943], expanded_key[944], expanded_key[945], expanded_key[946], expanded_key[947], expanded_key[948], expanded_key[949], expanded_key[950], expanded_key[951], expanded_key[952], expanded_key[953], expanded_key[954], expanded_key[955], expanded_key[956], expanded_key[957], expanded_key[958], expanded_key[959], expanded_key[960], expanded_key[961], expanded_key[962], expanded_key[963], expanded_key[964], expanded_key[965], expanded_key[966], expanded_key[967], expanded_key[968], expanded_key[969], expanded_key[970], expanded_key[971], expanded_key[972], expanded_key[973], expanded_key[974], expanded_key[975], expanded_key[976], expanded_key[977], expanded_key[978], expanded_key[979], expanded_key[980], expanded_key[981], expanded_key[982], expanded_key[983], expanded_key[984], expanded_key[985], expanded_key[986], expanded_key[987], expanded_key[988], expanded_key[989], expanded_key[990], expanded_key[991], expanded_key[992], expanded_key[993], expanded_key[994], expanded_key[995], expanded_key[996], expanded_key[997], expanded_key[998], expanded_key[999], expanded_key[1000], expanded_key[1001], expanded_key[1002], expanded_key[1003], expanded_key[1004], expanded_key[1005], expanded_key[1006], expanded_key[1007], expanded_key[1008], expanded_key[1009], expanded_key[1010], expanded_key[1011], expanded_key[1012], expanded_key[1013], expanded_key[1014], expanded_key[1015], expanded_key[1016], expanded_key[1017], expanded_key[1018], expanded_key[1019], expanded_key[1020], expanded_key[1021], expanded_key[1022], expanded_key[1023]};
    assign temp_11 = new_8;
    assign tmp1985 = tmp1983 ^ tmp1984;
    assign substituted_w23 = tmp150;
    assign tmp1129 = tmp1127 ^ tmp1128;
        assign tmp1325 = mem_7[tmp1258];
        assign tmp2288 = mem_6[tmp2181];
    assign tmp1041 = tmp1078;
    assign tmp1438 = {temp_21[72], temp_21[73], temp_21[74], temp_21[75], temp_21[76], temp_21[77], temp_21[78], temp_21[79]};
    assign tmp352 = tmp396;
    assign tmp623 = tmp621 ^ tmp622;
    assign c3_w23 = tmp148;
    assign tmp1070 = {tmp1069[0], tmp1069[1], tmp1069[2], tmp1069[3], tmp1069[4], tmp1069[5], tmp1069[6], tmp1069[7]};
    assign tmp63 = {tmp61[16], tmp61[17], tmp61[18], tmp61[19], tmp61[20], tmp61[21], tmp61[22], tmp61[23]};
    assign tmp37 = {tmp36[24], tmp36[25], tmp36[26], tmp36[27], tmp36[28], tmp36[29], tmp36[30], tmp36[31]};
    assign tmp587 = tmp666;
    assign tmp1228 = tmp1244;
    assign tmp1183 = tmp1184;
    assign tmp345 = {temp_3[24], temp_3[25], temp_3[26], temp_3[27], temp_3[28], temp_3[29], temp_3[30], temp_3[31]};
        assign tmp940 = mem_6[tmp805];
    assign tmp483 = tmp481 ^ tmp482;
        assign tmp1342 = mem_5[tmp1257];
    assign tmp2144 = tmp2160;
        assign tmp2208 = mem_6[tmp2175];
    assign tmp1562 = {tmp1561[0], tmp1561[1], tmp1561[2], tmp1561[3], tmp1561[4], tmp1561[5], tmp1561[6], tmp1561[7]};
    assign tmp2065 = tmp2063 ^ tmp2064;
    assign tmp569 = {temp_7[72], temp_7[73], temp_7[74], temp_7[75], temp_7[76], temp_7[77], temp_7[78], temp_7[79]};
    assign tmp1093 = tmp1091 ^ tmp1092;
        assign tmp1842 = mem_5[tmp1726];
    assign tmp208 = tmp183 ^ xor_w31;
        assign tmp422 = mem_5[tmp337];
    assign tmp1681 = tmp1697;
    assign tmp2375 = tmp2391;
        assign tmp1127 = mem_7[tmp1032];
    assign tmp1503 = tmp1554;
        assign tmp1112 = mem_5[tmp1027];
    assign tmp113 = {tmp111[16], tmp111[17], tmp111[18], tmp111[19], tmp111[20], tmp111[21], tmp111[22], tmp111[23]};
    assign tmp1667 = {temp_25[80], temp_25[81], temp_25[82], temp_25[83], temp_25[84], temp_25[85], temp_25[86], temp_25[87]};
        assign tmp418 = mem_4[tmp338];
    assign tmp2263 = tmp2261 ^ tmp2262;
    assign tmp714 = {tmp713[0], tmp713[1], tmp713[2], tmp713[3], tmp713[4], tmp713[5], tmp713[6], tmp713[7]};
    assign tmp260 = tmp259 ^ tmp235;
    assign tmp2078 = {tmp2077[0], tmp2077[1], tmp2077[2], tmp2077[3], tmp2077[4], tmp2077[5], tmp2077[6], tmp2077[7]};
    assign tmp1553 = tmp1551 ^ tmp1552;
    assign tmp572 = {temp_7[48], temp_7[49], temp_7[50], temp_7[51], temp_7[52], temp_7[53], temp_7[54], temp_7[55]};
    assign tmp1541 = tmp1539 ^ tmp1540;
        assign tmp21 = mem_1[b1_w3];
    assign tmp2094 = {tmp2093[0], tmp2093[1], tmp2093[2], tmp2093[3], tmp2093[4], tmp2093[5], tmp2093[6], tmp2093[7]};
    assign c1_w11 = tmp71;
    assign tmp1499 = tmp1522;
        assign tmp2298 = mem_4[tmp2183];
    assign substituted_w39 = tmp250;
    assign tmp2145 = tmp2161;
    assign tmp1896 = {temp_29[88], temp_29[89], temp_29[90], temp_29[91], temp_29[92], temp_29[93], temp_29[94], temp_29[95]};
    assign tmp526 = {temp_5[8], temp_5[9], temp_5[10], temp_5[11], temp_5[12], temp_5[13], temp_5[14], temp_5[15]};
    assign tmp1736 = tmp1808;
    assign tmp1979 = tmp1977 ^ tmp1978;
    assign a1_w31 = tmp187;
    assign tmp2019 = tmp2017 ^ tmp2018;
    assign tmp415 = tmp413 ^ tmp414;
        assign tmp1574 = mem_6[tmp1488];
        assign tmp890 = mem_5[tmp802];
    assign tmp713 = tmp711 ^ tmp712;
    assign tmp1678 = tmp1694;
    assign tmp607 = tmp605 ^ tmp606;
    assign c3_w7 = tmp48;
        assign tmp676 = mem_5[tmp574];
        assign tmp2156 = mem_2[tmp2124];
        assign tmp22 = mem_1[b2_w3];
    assign tmp735 = {temp_8[40], temp_8[41], temp_8[42], temp_8[43], temp_8[44], temp_8[45], temp_8[46], temp_8[47]};
    assign tmp86 = tmp85 ^ tmp61;
    assign tmp799 = {temp_11[72], temp_11[73], temp_11[74], temp_11[75], temp_11[76], temp_11[77], temp_11[78], temp_11[79]};
    assign tmp679 = tmp677 ^ tmp678;
    assign tmp1364 = {tmp1363[0], tmp1363[1], tmp1363[2], tmp1363[3], tmp1363[4], tmp1363[5], tmp1363[6], tmp1363[7]};
        assign tmp603 = mem_7[tmp564];
        assign tmp1702 = mem_2[tmp1670];
    assign tmp2365 = {temp_37[16], temp_37[17], temp_37[18], temp_37[19], temp_37[20], temp_37[21], temp_37[22], temp_37[23]};
    assign tmp759 = tmp775;
    assign tmp338 = {temp_3[80], temp_3[81], temp_3[82], temp_3[83], temp_3[84], temp_3[85], temp_3[86], temp_3[87]};
    assign temp_31 = new_3;
    assign tmp1957 = {temp_31[8], temp_31[9], temp_31[10], temp_31[11], temp_31[12], temp_31[13], temp_31[14], temp_31[15]};
    assign tmp2108 = {temp_32[96], temp_32[97], temp_32[98], temp_32[99], temp_32[100], temp_32[101], temp_32[102], temp_32[103]};
        assign tmp1176 = mem_5[tmp1035];
    assign tmp1797 = tmp1795 ^ tmp1796;
        assign tmp2072 = mem_5[tmp1956];
        assign tmp52 = mem_3[const51_2];
    assign concat_w11 = tmp81;
    assign tmp1078 = {tmp1077[0], tmp1077[1], tmp1077[2], tmp1077[3], tmp1077[4], tmp1077[5], tmp1077[6], tmp1077[7]};
    assign tmp1444 = {temp_21[24], temp_21[25], temp_21[26], temp_21[27], temp_21[28], temp_21[29], temp_21[30], temp_21[31]};
    assign tmp772 = tmp788;
        assign tmp1237 = mem_2[tmp1205];
    assign tmp2099 = tmp2097 ^ tmp2098;
        assign tmp844 = mem_6[tmp793];
    assign tmp1121 = tmp1119 ^ tmp1120;
        assign tmp1750 = mem_4[tmp1716];
        assign tmp557 = mem_2[tmp525];
    assign tmp634 = {tmp633[0], tmp633[1], tmp633[2], tmp633[3], tmp633[4], tmp633[5], tmp633[6], tmp633[7]};
        assign tmp2261 = mem_7[tmp2180];
        assign tmp2274 = mem_4[tmp2184];
    assign tmp1369 = tmp1367 ^ tmp1368;
        assign tmp1344 = mem_6[tmp1258];
        assign tmp2206 = mem_5[tmp2174];
    assign tmp1022 = temp_14 ^ tmp1021;
        assign tmp1285 = mem_7[tmp1253];
    assign tmp340 = {temp_3[64], temp_3[65], temp_3[66], temp_3[67], temp_3[68], temp_3[69], temp_3[70], temp_3[71]};
        assign tmp386 = mem_4[tmp334];
    assign tmp1023 = {temp_15[120], temp_15[121], temp_15[122], temp_15[123], temp_15[124], temp_15[125], temp_15[126], temp_15[127]};
        assign tmp1836 = mem_6[tmp1722];
        assign tmp1245 = mem_2[tmp1213];
    assign tmp2124 = {temp_33[104], temp_33[105], temp_33[106], temp_33[107], temp_33[108], temp_33[109], temp_33[110], temp_33[111]};
        assign tmp1394 = mem_4[tmp1265];
        assign tmp2066 = mem_6[tmp1952];
        assign tmp1156 = mem_4[tmp1038];
    assign tmp955 = {temp_12[120], temp_12[121], temp_12[122], temp_12[123], temp_12[124], temp_12[125], temp_12[126], temp_12[127]};
        assign tmp2032 = mem_5[tmp1947];
    assign tmp311 = tmp327;
        assign tmp46 = mem_1[b1_w7];
        assign tmp2306 = mem_4[tmp2188];
    assign tmp797 = {temp_11[88], temp_11[89], temp_11[90], temp_11[91], temp_11[92], temp_11[93], temp_11[94], temp_11[95]};
    assign tmp2198 = tmp2284;
    assign tmp272 = {new_state[64], new_state[65], new_state[66], new_state[67], new_state[68], new_state[69], new_state[70], new_state[71]};
    assign tmp2203 = tmp2324;
    assign tmp1094 = {tmp1093[0], tmp1093[1], tmp1093[2], tmp1093[3], tmp1093[4], tmp1093[5], tmp1093[6], tmp1093[7]};
        assign tmp1235 = mem_2[tmp1203];
        assign tmp1588 = mem_5[tmp1493];
        assign tmp1785 = mem_7[tmp1718];
    assign tmp1409 = tmp1407 ^ tmp1408;
        assign tmp1852 = mem_6[tmp1728];
        assign tmp314 = mem_2[tmp282];
        assign tmp1018 = mem_2[tmp986];
    assign tmp269 = {new_state[88], new_state[89], new_state[90], new_state[91], new_state[92], new_state[93], new_state[94], new_state[95]};
    assign tmp34 = tmp33 ^ tmp9;
        assign tmp461 = mem_7[tmp345];
        assign tmp1818 = mem_5[tmp1723];
    assign tmp681 = tmp679 ^ tmp680;
        assign tmp948 = mem_6[tmp806];
        assign tmp1368 = mem_6[tmp1261];
        assign tmp716 = mem_5[tmp575];
    assign tmp594 = tmp722;
        assign tmp1373 = mem_7[tmp1264];
        assign tmp1408 = mem_6[tmp1266];
    assign tmp2093 = tmp2091 ^ tmp2092;
        assign tmp224 = mem_1[b4_w35];
    assign tmp447 = tmp445 ^ tmp446;
    assign tmp145 = {shifted_w23[0], shifted_w23[1], shifted_w23[2], shifted_w23[3], shifted_w23[4], shifted_w23[5], shifted_w23[6], shifted_w23[7]};
    assign tmp1407 = tmp1405 ^ tmp1406;
    assign tmp839 = tmp837 ^ tmp838;
    assign tmp739 = {temp_8[8], temp_8[9], temp_8[10], temp_8[11], temp_8[12], temp_8[13], temp_8[14], temp_8[15]};
        assign tmp1242 = mem_2[tmp1210];
    assign tmp2143 = tmp2159;
        assign tmp2031 = mem_7[tmp1950];
        assign tmp2056 = mem_5[tmp1954];
    assign rc4_w27 = const180_0;
    assign tmp2062 = {tmp2061[0], tmp2061[1], tmp2061[2], tmp2061[3], tmp2061[4], tmp2061[5], tmp2061[6], tmp2061[7]};
        assign tmp2326 = mem_5[tmp2185];
    assign tmp494 = {tmp349, tmp350, tmp351, tmp352, tmp353, tmp354, tmp355, tmp356, tmp357, tmp358, tmp359, tmp360, tmp361, tmp362, tmp363, tmp364};
    assign tmp243 = {shifted_w39[16], shifted_w39[17], shifted_w39[18], shifted_w39[19], shifted_w39[20], shifted_w39[21], shifted_w39[22], shifted_w39[23]};
        assign tmp2210 = mem_4[tmp2176];
    assign new_2 = tmp2172;
    assign tmp1521 = tmp1519 ^ tmp1520;
        assign tmp2394 = mem_2[tmp2362];
    assign tmp59 = tmp58 ^ tmp34;
    assign tmp2117 = {temp_32[24], temp_32[25], temp_32[26], temp_32[27], temp_32[28], temp_32[29], temp_32[30], temp_32[31]};
    assign tmp1672 = {temp_25[40], temp_25[41], temp_25[42], temp_25[43], temp_25[44], temp_25[45], temp_25[46], temp_25[47]};
    assign b2_w23 = tmp143;
    assign rc2_w35 = const228_0;
        assign tmp1640 = mem_4[tmp1497];
        assign tmp1475 = mem_2[tmp1443];
        assign tmp2100 = mem_4[tmp1957];
        assign tmp121 = mem_1[b1_w19];
    assign tmp1511 = tmp1618;
    assign tmp2196 = tmp2268;
    assign tmp245 = {shifted_w39[0], shifted_w39[1], shifted_w39[2], shifted_w39[3], shifted_w39[4], shifted_w39[5], shifted_w39[6], shifted_w39[7]};
    assign tmp210 = tmp209 ^ tmp185;
    assign tmp1215 = {temp_17[16], temp_17[17], temp_17[18], temp_17[19], temp_17[20], temp_17[21], temp_17[22], temp_17[23]};
    assign tmp962 = {temp_12[64], temp_12[65], temp_12[66], temp_12[67], temp_12[68], temp_12[69], temp_12[70], temp_12[71]};
        assign tmp1164 = mem_4[tmp1035];
    assign tmp2307 = tmp2305 ^ tmp2306;
    assign c2_w35 = tmp222;
        assign tmp1793 = mem_7[tmp1719];
    assign tmp354 = tmp412;
    assign tmp372 = {tmp371[0], tmp371[1], tmp371[2], tmp371[3], tmp371[4], tmp371[5], tmp371[6], tmp371[7]};
        assign tmp1148 = mem_4[tmp1033];
    assign tmp436 = {tmp435[0], tmp435[1], tmp435[2], tmp435[3], tmp435[4], tmp435[5], tmp435[6], tmp435[7]};
    assign tmp1906 = {temp_29[8], temp_29[9], temp_29[10], temp_29[11], temp_29[12], temp_29[13], temp_29[14], temp_29[15]};
        assign tmp2048 = mem_5[tmp1953];
    assign tmp2041 = tmp2039 ^ tmp2040;
    assign tmp2153 = tmp2169;
        assign tmp1622 = mem_6[tmp1498];
        assign tmp2008 = mem_5[tmp1948];
    assign tmp336 = {temp_3[96], temp_3[97], temp_3[98], temp_3[99], temp_3[100], temp_3[101], temp_3[102], temp_3[103]};
        assign tmp424 = mem_6[tmp338];
        assign tmp147 = mem_1[b2_w23];
    assign tmp1186 = {temp_16[112], temp_16[113], temp_16[114], temp_16[115], temp_16[116], temp_16[117], temp_16[118], temp_16[119]};
        assign tmp1306 = mem_4[tmp1254];
    assign rc4_w23 = const155_0;
    assign tmp2291 = tmp2289 ^ tmp2290;
    assign tmp2363 = {temp_37[32], temp_37[33], temp_37[34], temp_37[35], temp_37[36], temp_37[37], temp_37[38], temp_37[39]};
    assign tmp1734 = tmp1792;
        assign tmp1746 = mem_5[tmp1714];
    assign tmp119 = {shifted_w19[8], shifted_w19[9], shifted_w19[10], shifted_w19[11], shifted_w19[12], shifted_w19[13], shifted_w19[14], shifted_w19[15]};
    assign tmp951 = tmp949 ^ tmp950;
    assign c2_w3 = tmp22;
    assign tmp8 = {aes_key[96], aes_key[97], aes_key[98], aes_key[99], aes_key[100], aes_key[101], aes_key[102], aes_key[103], aes_key[104], aes_key[105], aes_key[106], aes_key[107], aes_key[108], aes_key[109], aes_key[110], aes_key[111], aes_key[112], aes_key[113], aes_key[114], aes_key[115], aes_key[116], aes_key[117], aes_key[118], aes_key[119], aes_key[120], aes_key[121], aes_key[122], aes_key[123], aes_key[124], aes_key[125], aes_key[126], aes_key[127]};
    assign b2_w19 = tmp118;
        assign tmp2010 = mem_6[tmp1949];
    assign tmp752 = {temp_9[40], temp_9[41], temp_9[42], temp_9[43], temp_9[44], temp_9[45], temp_9[46], temp_9[47]};
        assign tmp720 = mem_4[tmp577];
    assign tmp581 = tmp618;
    assign tmp220 = {shifted_w35[0], shifted_w35[1], shifted_w35[2], shifted_w35[3], shifted_w35[4], shifted_w35[5], shifted_w35[6], shifted_w35[7]};
        assign tmp1825 = mem_7[tmp1723];
    assign tmp332 = temp_2 ^ tmp331;
    assign tmp896 = {tmp895[0], tmp895[1], tmp895[2], tmp895[3], tmp895[4], tmp895[5], tmp895[6], tmp895[7]};
        assign tmp2317 = mem_7[tmp2187];
    assign tmp2308 = {tmp2307[0], tmp2307[1], tmp2307[2], tmp2307[3], tmp2307[4], tmp2307[5], tmp2307[6], tmp2307[7]};
    assign c3_w31 = tmp198;
    assign tmp563 = {temp_7[120], temp_7[121], temp_7[122], temp_7[123], temp_7[124], temp_7[125], temp_7[126], temp_7[127]};
    assign tmp762 = tmp778;
        assign tmp325 = mem_2[tmp293];
    assign tmp301 = tmp317;
    assign tmp1874 = {tmp1729, tmp1730, tmp1731, tmp1732, tmp1733, tmp1734, tmp1735, tmp1736, tmp1737, tmp1738, tmp1739, tmp1740, tmp1741, tmp1742, tmp1743, tmp1744};
        assign tmp1016 = mem_2[tmp984];
    assign tmp527 = {temp_5[0], temp_5[1], temp_5[2], temp_5[3], temp_5[4], temp_5[5], temp_5[6], temp_5[7]};
    assign tmp1829 = tmp1827 ^ tmp1828;
    assign tmp169 = {shifted_w27[8], shifted_w27[9], shifted_w27[10], shifted_w27[11], shifted_w27[12], shifted_w27[13], shifted_w27[14], shifted_w27[15]};
        assign tmp1066 = mem_6[tmp1026];
        assign tmp1994 = mem_6[tmp1943];
    assign tmp771 = tmp787;
    assign tmp1198 = {temp_16[16], temp_16[17], temp_16[18], temp_16[19], temp_16[20], temp_16[21], temp_16[22], temp_16[23]};
    assign a2_w27 = tmp163;
    assign tmp138 = {tmp136[16], tmp136[17], tmp136[18], tmp136[19], tmp136[20], tmp136[21], tmp136[22], tmp136[23]};
        assign tmp1336 = mem_6[tmp1257];
    assign tmp2319 = tmp2317 ^ tmp2318;
    assign tmp1643 = tmp1644;
    assign tmp289 = {temp_1[64], temp_1[65], temp_1[66], temp_1[67], temp_1[68], temp_1[69], temp_1[70], temp_1[71]};
    assign tmp1912 = tmp1928;
    assign rc2_w31 = const203_0;
    assign tmp1652 = {temp_24[64], temp_24[65], temp_24[66], temp_24[67], temp_24[68], temp_24[69], temp_24[70], temp_24[71]};
    assign tmp2327 = tmp2325 ^ tmp2326;
    assign tmp403 = tmp401 ^ tmp402;
    assign tmp1773 = tmp1771 ^ tmp1772;
        assign tmp485 = mem_7[tmp348];
    assign tmp2350 = {temp_36[0], temp_36[1], temp_36[2], temp_36[3], temp_36[4], temp_36[5], temp_36[6], temp_36[7]};
    assign tmp491 = tmp489 ^ tmp490;
        assign tmp324 = mem_2[tmp292];
    assign tmp1363 = tmp1361 ^ tmp1362;
    assign tmp645 = tmp643 ^ tmp644;
        assign tmp474 = mem_4[tmp345];
    assign tmp1731 = tmp1768;
    assign tmp214 = {tmp211[8], tmp211[9], tmp211[10], tmp211[11], tmp211[12], tmp211[13], tmp211[14], tmp211[15]};
    assign tmp693 = tmp691 ^ tmp692;
    assign tmp1958 = {temp_31[0], temp_31[1], temp_31[2], temp_31[3], temp_31[4], temp_31[5], temp_31[6], temp_31[7]};
    assign tmp1626 = {tmp1625[0], tmp1625[1], tmp1625[2], tmp1625[3], tmp1625[4], tmp1625[5], tmp1625[6], tmp1625[7]};
    assign a1_w19 = tmp112;
    assign tmp2109 = {temp_32[88], temp_32[89], temp_32[90], temp_32[91], temp_32[92], temp_32[93], temp_32[94], temp_32[95]};
    assign tmp845 = tmp843 ^ tmp844;
    assign tmp626 = {tmp625[0], tmp625[1], tmp625[2], tmp625[3], tmp625[4], tmp625[5], tmp625[6], tmp625[7]};
    assign tmp971 = {tmp955, tmp968, tmp965, tmp962, tmp959, tmp956, tmp969, tmp966, tmp963, tmp960, tmp957, tmp970, tmp967, tmp964, tmp961, tmp958};
    assign tmp1631 = tmp1629 ^ tmp1630;
    assign tmp1037 = {temp_15[8], temp_15[9], temp_15[10], temp_15[11], temp_15[12], temp_15[13], temp_15[14], temp_15[15]};
    assign tmp2053 = tmp2051 ^ tmp2052;
    assign tmp859 = tmp857 ^ tmp858;
        assign tmp2076 = mem_4[tmp1958];
    assign tmp2176 = {temp_35[96], temp_35[97], temp_35[98], temp_35[99], temp_35[100], temp_35[101], temp_35[102], temp_35[103]};
        assign tmp1844 = mem_6[tmp1727];
        assign tmp49 = mem_1[b4_w7];
    assign tmp2104 = {tmp1959, tmp1960, tmp1961, tmp1962, tmp1963, tmp1964, tmp1965, tmp1966, tmp1967, tmp1968, tmp1969, tmp1970, tmp1971, tmp1972, tmp1973, tmp1974};
    assign tmp502 = {temp_4[64], temp_4[65], temp_4[66], temp_4[67], temp_4[68], temp_4[69], temp_4[70], temp_4[71]};
    assign tmp847 = tmp845 ^ tmp846;
    assign tmp505 = {temp_4[40], temp_4[41], temp_4[42], temp_4[43], temp_4[44], temp_4[45], temp_4[46], temp_4[47]};
        assign tmp48 = mem_1[b3_w7];
    assign tmp2067 = tmp2065 ^ tmp2066;
    assign c4_w7 = tmp49;
        assign tmp1095 = mem_7[tmp1028];
    assign tmp2030 = {tmp2029[0], tmp2029[1], tmp2029[2], tmp2029[3], tmp2029[4], tmp2029[5], tmp2029[6], tmp2029[7]};
    assign tmp346 = {temp_3[16], temp_3[17], temp_3[18], temp_3[19], temp_3[20], temp_3[21], temp_3[22], temp_3[23]};
    assign input_wire_6 = temp_18;
        assign tmp1072 = mem_5[tmp1026];
    assign c4_w27 = tmp174;
    assign tmp191 = {a2_w31, a3_w31, a4_w31, a1_w31};
    assign tmp1404 = {tmp1403[0], tmp1403[1], tmp1403[2], tmp1403[3], tmp1403[4], tmp1403[5], tmp1403[6], tmp1403[7]};
    assign tmp998 = tmp1014;
    assign tmp1038 = {temp_15[0], temp_15[1], temp_15[2], temp_15[3], temp_15[4], temp_15[5], temp_15[6], temp_15[7]};
    assign tmp1263 = {temp_19[40], temp_19[41], temp_19[42], temp_19[43], temp_19[44], temp_19[45], temp_19[46], temp_19[47]};
    assign tmp1909 = tmp1925;
    assign tmp2190 = tmp2220;
        assign tmp74 = mem_1[b4_w11];
    assign tmp313 = tmp329;
    assign tmp861 = tmp859 ^ tmp860;
        assign tmp1471 = mem_2[tmp1439];
    assign tmp809 = tmp832;
    assign a2_w35 = tmp213;
        assign tmp2068 = mem_4[tmp1953];
    assign tmp1671 = {temp_25[48], temp_25[49], temp_25[50], temp_25[51], temp_25[52], temp_25[53], temp_25[54], temp_25[55]};
    assign tmp747 = {temp_9[80], temp_9[81], temp_9[82], temp_9[83], temp_9[84], temp_9[85], temp_9[86], temp_9[87]};
        assign tmp1473 = mem_2[tmp1441];
    assign tmp520 = {temp_5[56], temp_5[57], temp_5[58], temp_5[59], temp_5[60], temp_5[61], temp_5[62], temp_5[63]};
        assign tmp1846 = mem_4[tmp1728];
        assign tmp1236 = mem_2[tmp1204];
    assign tmp1839 = tmp1837 ^ tmp1838;
    assign tmp1659 = {temp_24[8], temp_24[9], temp_24[10], temp_24[11], temp_24[12], temp_24[13], temp_24[14], temp_24[15]};
    assign tmp703 = tmp701 ^ tmp702;
    assign tmp2367 = {temp_37[0], temp_37[1], temp_37[2], temp_37[3], temp_37[4], temp_37[5], temp_37[6], temp_37[7]};
    assign tmp2130 = {temp_33[56], temp_33[57], temp_33[58], temp_33[59], temp_33[60], temp_33[61], temp_33[62], temp_33[63]};
    assign tmp695 = tmp693 ^ tmp694;
    assign tmp1719 = {temp_27[72], temp_27[73], temp_27[74], temp_27[75], temp_27[76], temp_27[77], temp_27[78], temp_27[79]};
    assign tmp2149 = tmp2165;
        assign tmp789 = mem_2[tmp757];
        assign tmp490 = mem_4[tmp347];
    assign tmp2324 = {tmp2323[0], tmp2323[1], tmp2323[2], tmp2323[3], tmp2323[4], tmp2323[5], tmp2323[6], tmp2323[7]};
        assign tmp2294 = mem_5[tmp2181];
    assign tmp2013 = tmp2011 ^ tmp2012;
        assign tmp916 = mem_6[tmp802];
    assign tmp2120 = {temp_32[0], temp_32[1], temp_32[2], temp_32[3], temp_32[4], temp_32[5], temp_32[6], temp_32[7]};
    assign tmp562 = temp_6 ^ tmp561;
    assign tmp242 = {shifted_w39[24], shifted_w39[25], shifted_w39[26], shifted_w39[27], shifted_w39[28], shifted_w39[29], shifted_w39[30], shifted_w39[31]};
    assign tmp2378 = tmp2394;
    assign tmp1668 = {temp_25[72], temp_25[73], temp_25[74], temp_25[75], temp_25[76], temp_25[77], temp_25[78], temp_25[79]};
        assign tmp1862 = mem_4[tmp1726];
        assign tmp1352 = mem_6[tmp1263];
    assign tmp748 = {temp_9[72], temp_9[73], temp_9[74], temp_9[75], temp_9[76], temp_9[77], temp_9[78], temp_9[79]};
    assign tmp369 = tmp367 ^ tmp368;
        assign tmp1341 = mem_7[tmp1260];
    assign tmp1377 = tmp1375 ^ tmp1376;
        assign tmp2253 = mem_7[tmp2179];
        assign tmp2385 = mem_2[tmp2353];
    assign tmp1962 = tmp2006;
        assign tmp390 = mem_5[tmp333];
    assign tmp1683 = tmp1699;
    assign tmp1949 = {temp_31[72], temp_31[73], temp_31[74], temp_31[75], temp_31[76], temp_31[77], temp_31[78], temp_31[79]};
    assign rc1_w23 = tmp152;
        assign tmp775 = mem_2[tmp743];
        assign tmp1572 = mem_5[tmp1487];
    assign tmp85 = tmp84 ^ tmp60;
    assign xor_w23 = tmp157;
    assign tmp931 = tmp929 ^ tmp930;
    assign tmp1021 = {expanded_key[512], expanded_key[513], expanded_key[514], expanded_key[515], expanded_key[516], expanded_key[517], expanded_key[518], expanded_key[519], expanded_key[520], expanded_key[521], expanded_key[522], expanded_key[523], expanded_key[524], expanded_key[525], expanded_key[526], expanded_key[527], expanded_key[528], expanded_key[529], expanded_key[530], expanded_key[531], expanded_key[532], expanded_key[533], expanded_key[534], expanded_key[535], expanded_key[536], expanded_key[537], expanded_key[538], expanded_key[539], expanded_key[540], expanded_key[541], expanded_key[542], expanded_key[543], expanded_key[544], expanded_key[545], expanded_key[546], expanded_key[547], expanded_key[548], expanded_key[549], expanded_key[550], expanded_key[551], expanded_key[552], expanded_key[553], expanded_key[554], expanded_key[555], expanded_key[556], expanded_key[557], expanded_key[558], expanded_key[559], expanded_key[560], expanded_key[561], expanded_key[562], expanded_key[563], expanded_key[564], expanded_key[565], expanded_key[566], expanded_key[567], expanded_key[568], expanded_key[569], expanded_key[570], expanded_key[571], expanded_key[572], expanded_key[573], expanded_key[574], expanded_key[575], expanded_key[576], expanded_key[577], expanded_key[578], expanded_key[579], expanded_key[580], expanded_key[581], expanded_key[582], expanded_key[583], expanded_key[584], expanded_key[585], expanded_key[586], expanded_key[587], expanded_key[588], expanded_key[589], expanded_key[590], expanded_key[591], expanded_key[592], expanded_key[593], expanded_key[594], expanded_key[595], expanded_key[596], expanded_key[597], expanded_key[598], expanded_key[599], expanded_key[600], expanded_key[601], expanded_key[602], expanded_key[603], expanded_key[604], expanded_key[605], expanded_key[606], expanded_key[607], expanded_key[608], expanded_key[609], expanded_key[610], expanded_key[611], expanded_key[612], expanded_key[613], expanded_key[614], expanded_key[615], expanded_key[616], expanded_key[617], expanded_key[618], expanded_key[619], expanded_key[620], expanded_key[621], expanded_key[622], expanded_key[623], expanded_key[624], expanded_key[625], expanded_key[626], expanded_key[627], expanded_key[628], expanded_key[629], expanded_key[630], expanded_key[631], expanded_key[632], expanded_key[633], expanded_key[634], expanded_key[635], expanded_key[636], expanded_key[637], expanded_key[638], expanded_key[639]};
    assign tmp1821 = tmp1819 ^ tmp1820;
    assign tmp441 = tmp439 ^ tmp440;
        assign tmp1080 = mem_5[tmp1023];
    assign tmp1182 = {tmp1181[0], tmp1181[1], tmp1181[2], tmp1181[3], tmp1181[4], tmp1181[5], tmp1181[6], tmp1181[7]};
    assign tmp831 = tmp829 ^ tmp830;
    assign tmp840 = {tmp839[0], tmp839[1], tmp839[2], tmp839[3], tmp839[4], tmp839[5], tmp839[6], tmp839[7]};
    assign tmp639 = tmp637 ^ tmp638;
    assign tmp353 = tmp404;
        assign tmp127 = mem_3[const126_5];
    assign tmp2267 = tmp2265 ^ tmp2266;
        assign tmp99 = mem_1[b4_w15];
    assign tmp375 = tmp373 ^ tmp374;
        assign tmp646 = mem_6[tmp567];
        assign tmp1160 = mem_5[tmp1037];
    assign tmp2243 = tmp2241 ^ tmp2242;
    assign tmp1873 = tmp1874;
    assign xor_w19 = tmp132;
    assign tmp685 = tmp683 ^ tmp684;
    assign tmp1546 = {tmp1545[0], tmp1545[1], tmp1545[2], tmp1545[3], tmp1545[4], tmp1545[5], tmp1545[6], tmp1545[7]};
    assign tmp1319 = tmp1317 ^ tmp1318;
    assign tmp1145 = tmp1143 ^ tmp1144;
        assign tmp612 = mem_5[tmp566];
    assign tmp207 = concat_w31 ^ substituted_w31;
    assign tmp1740 = tmp1840;
    assign tmp2339 = {temp_36[88], temp_36[89], temp_36[90], temp_36[91], temp_36[92], temp_36[93], temp_36[94], temp_36[95]};
    assign c4_w3 = tmp24;
        assign tmp926 = mem_4[tmp808];
        assign tmp1542 = mem_6[tmp1484];
    assign tmp724 = {tmp579, tmp580, tmp581, tmp582, tmp583, tmp584, tmp585, tmp586, tmp587, tmp588, tmp589, tmp590, tmp591, tmp592, tmp593, tmp594};
    assign tmp2181 = {temp_35[56], temp_35[57], temp_35[58], temp_35[59], temp_35[60], temp_35[61], temp_35[62], temp_35[63]};
    assign tmp1048 = tmp1134;
        assign tmp945 = mem_7[tmp808];
        assign tmp172 = mem_1[b2_w27];
    assign tmp1383 = tmp1381 ^ tmp1382;
    assign tmp773 = tmp789;
        assign tmp2390 = mem_2[tmp2358];
    assign tmp1351 = tmp1349 ^ tmp1350;
        assign tmp559 = mem_2[tmp527];
    assign tmp528 = tmp544;
    assign rc2_w3 = const28_0;
    assign xor_w35 = tmp232;
    assign tmp1379 = tmp1377 ^ tmp1378;
    assign tmp534 = tmp550;
        assign tmp876 = mem_6[tmp797];
    assign tmp380 = {tmp379[0], tmp379[1], tmp379[2], tmp379[3], tmp379[4], tmp379[5], tmp379[6], tmp379[7]};
    assign tmp719 = tmp717 ^ tmp718;
        assign tmp1296 = mem_6[tmp1256];
    assign tmp811 = tmp848;
    assign tmp1755 = tmp1753 ^ tmp1754;
    assign rc1_w35 = tmp227;
    assign tmp68 = {shifted_w11[16], shifted_w11[17], shifted_w11[18], shifted_w11[19], shifted_w11[20], shifted_w11[21], shifted_w11[22], shifted_w11[23]};
    assign tmp84 = tmp83 ^ tmp59;
    assign tmp218 = {shifted_w35[16], shifted_w35[17], shifted_w35[18], shifted_w35[19], shifted_w35[20], shifted_w35[21], shifted_w35[22], shifted_w35[23]};
    assign tmp982 = {temp_13[40], temp_13[41], temp_13[42], temp_13[43], temp_13[44], temp_13[45], temp_13[46], temp_13[47]};
    assign tmp134 = tmp133 ^ tmp109;
    assign tmp2171 = {expanded_key[1152], expanded_key[1153], expanded_key[1154], expanded_key[1155], expanded_key[1156], expanded_key[1157], expanded_key[1158], expanded_key[1159], expanded_key[1160], expanded_key[1161], expanded_key[1162], expanded_key[1163], expanded_key[1164], expanded_key[1165], expanded_key[1166], expanded_key[1167], expanded_key[1168], expanded_key[1169], expanded_key[1170], expanded_key[1171], expanded_key[1172], expanded_key[1173], expanded_key[1174], expanded_key[1175], expanded_key[1176], expanded_key[1177], expanded_key[1178], expanded_key[1179], expanded_key[1180], expanded_key[1181], expanded_key[1182], expanded_key[1183], expanded_key[1184], expanded_key[1185], expanded_key[1186], expanded_key[1187], expanded_key[1188], expanded_key[1189], expanded_key[1190], expanded_key[1191], expanded_key[1192], expanded_key[1193], expanded_key[1194], expanded_key[1195], expanded_key[1196], expanded_key[1197], expanded_key[1198], expanded_key[1199], expanded_key[1200], expanded_key[1201], expanded_key[1202], expanded_key[1203], expanded_key[1204], expanded_key[1205], expanded_key[1206], expanded_key[1207], expanded_key[1208], expanded_key[1209], expanded_key[1210], expanded_key[1211], expanded_key[1212], expanded_key[1213], expanded_key[1214], expanded_key[1215], expanded_key[1216], expanded_key[1217], expanded_key[1218], expanded_key[1219], expanded_key[1220], expanded_key[1221], expanded_key[1222], expanded_key[1223], expanded_key[1224], expanded_key[1225], expanded_key[1226], expanded_key[1227], expanded_key[1228], expanded_key[1229], expanded_key[1230], expanded_key[1231], expanded_key[1232], expanded_key[1233], expanded_key[1234], expanded_key[1235], expanded_key[1236], expanded_key[1237], expanded_key[1238], expanded_key[1239], expanded_key[1240], expanded_key[1241], expanded_key[1242], expanded_key[1243], expanded_key[1244], expanded_key[1245], expanded_key[1246], expanded_key[1247], expanded_key[1248], expanded_key[1249], expanded_key[1250], expanded_key[1251], expanded_key[1252], expanded_key[1253], expanded_key[1254], expanded_key[1255], expanded_key[1256], expanded_key[1257], expanded_key[1258], expanded_key[1259], expanded_key[1260], expanded_key[1261], expanded_key[1262], expanded_key[1263], expanded_key[1264], expanded_key[1265], expanded_key[1266], expanded_key[1267], expanded_key[1268], expanded_key[1269], expanded_key[1270], expanded_key[1271], expanded_key[1272], expanded_key[1273], expanded_key[1274], expanded_key[1275], expanded_key[1276], expanded_key[1277], expanded_key[1278], expanded_key[1279]};
        assign tmp1616 = mem_4[tmp1498];
        assign tmp1159 = mem_7[tmp1036];
    assign tmp2241 = tmp2239 ^ tmp2240;
    assign tmp41 = {a2_w7, a3_w7, a4_w7, a1_w7};
    assign tmp2228 = {tmp2227[0], tmp2227[1], tmp2227[2], tmp2227[3], tmp2227[4], tmp2227[5], tmp2227[6], tmp2227[7]};
        assign tmp73 = mem_1[b3_w11];
    assign rc4_w19 = const130_0;
    assign tmp1040 = tmp1070;
        assign tmp548 = mem_2[tmp516];
    assign tmp661 = tmp659 ^ tmp660;
    assign tmp435 = tmp433 ^ tmp434;
    assign tmp1454 = tmp1470;
        assign tmp2232 = mem_6[tmp2174];
    assign tmp396 = {tmp395[0], tmp395[1], tmp395[2], tmp395[3], tmp395[4], tmp395[5], tmp395[6], tmp395[7]};
        assign tmp389 = mem_7[tmp336];
    assign tmp1188 = {temp_16[96], temp_16[97], temp_16[98], temp_16[99], temp_16[100], temp_16[101], temp_16[102], temp_16[103]};
    assign tmp304 = tmp320;
        assign tmp24 = mem_1[b4_w3];
    assign tmp333 = {temp_3[120], temp_3[121], temp_3[122], temp_3[123], temp_3[124], temp_3[125], temp_3[126], temp_3[127]};
        assign tmp102 = mem_3[const101_4];
    assign tmp268 = {new_state[96], new_state[97], new_state[98], new_state[99], new_state[100], new_state[101], new_state[102], new_state[103]};
        assign tmp857 = mem_7[tmp797];
    assign tmp988 = tmp1004;
    assign tmp1380 = {tmp1379[0], tmp1379[1], tmp1379[2], tmp1379[3], tmp1379[4], tmp1379[5], tmp1379[6], tmp1379[7]};
    assign tmp1889 = {temp_28[8], temp_28[9], temp_28[10], temp_28[11], temp_28[12], temp_28[13], temp_28[14], temp_28[15]};
    assign tmp1039 = tmp1062;
    assign tmp288 = {temp_1[72], temp_1[73], temp_1[74], temp_1[75], temp_1[76], temp_1[77], temp_1[78], temp_1[79]};
    assign rc2_w19 = const128_0;
    assign tmp1510 = tmp1610;
    assign tmp1664 = {temp_25[104], temp_25[105], temp_25[106], temp_25[107], temp_25[108], temp_25[109], temp_25[110], temp_25[111]};
    assign tmp1000 = tmp1016;
    assign tmp1085 = tmp1083 ^ tmp1084;
    assign tmp1625 = tmp1623 ^ tmp1624;
    assign tmp2382 = tmp2398;
    assign tmp1941 = {expanded_key[1024], expanded_key[1025], expanded_key[1026], expanded_key[1027], expanded_key[1028], expanded_key[1029], expanded_key[1030], expanded_key[1031], expanded_key[1032], expanded_key[1033], expanded_key[1034], expanded_key[1035], expanded_key[1036], expanded_key[1037], expanded_key[1038], expanded_key[1039], expanded_key[1040], expanded_key[1041], expanded_key[1042], expanded_key[1043], expanded_key[1044], expanded_key[1045], expanded_key[1046], expanded_key[1047], expanded_key[1048], expanded_key[1049], expanded_key[1050], expanded_key[1051], expanded_key[1052], expanded_key[1053], expanded_key[1054], expanded_key[1055], expanded_key[1056], expanded_key[1057], expanded_key[1058], expanded_key[1059], expanded_key[1060], expanded_key[1061], expanded_key[1062], expanded_key[1063], expanded_key[1064], expanded_key[1065], expanded_key[1066], expanded_key[1067], expanded_key[1068], expanded_key[1069], expanded_key[1070], expanded_key[1071], expanded_key[1072], expanded_key[1073], expanded_key[1074], expanded_key[1075], expanded_key[1076], expanded_key[1077], expanded_key[1078], expanded_key[1079], expanded_key[1080], expanded_key[1081], expanded_key[1082], expanded_key[1083], expanded_key[1084], expanded_key[1085], expanded_key[1086], expanded_key[1087], expanded_key[1088], expanded_key[1089], expanded_key[1090], expanded_key[1091], expanded_key[1092], expanded_key[1093], expanded_key[1094], expanded_key[1095], expanded_key[1096], expanded_key[1097], expanded_key[1098], expanded_key[1099], expanded_key[1100], expanded_key[1101], expanded_key[1102], expanded_key[1103], expanded_key[1104], expanded_key[1105], expanded_key[1106], expanded_key[1107], expanded_key[1108], expanded_key[1109], expanded_key[1110], expanded_key[1111], expanded_key[1112], expanded_key[1113], expanded_key[1114], expanded_key[1115], expanded_key[1116], expanded_key[1117], expanded_key[1118], expanded_key[1119], expanded_key[1120], expanded_key[1121], expanded_key[1122], expanded_key[1123], expanded_key[1124], expanded_key[1125], expanded_key[1126], expanded_key[1127], expanded_key[1128], expanded_key[1129], expanded_key[1130], expanded_key[1131], expanded_key[1132], expanded_key[1133], expanded_key[1134], expanded_key[1135], expanded_key[1136], expanded_key[1137], expanded_key[1138], expanded_key[1139], expanded_key[1140], expanded_key[1141], expanded_key[1142], expanded_key[1143], expanded_key[1144], expanded_key[1145], expanded_key[1146], expanded_key[1147], expanded_key[1148], expanded_key[1149], expanded_key[1150], expanded_key[1151]};
    assign tmp2192 = tmp2236;
    assign xor_w3 = tmp32;
    assign tmp741 = {tmp725, tmp738, tmp735, tmp732, tmp729, tmp726, tmp739, tmp736, tmp733, tmp730, tmp727, tmp740, tmp737, tmp734, tmp731, tmp728};
    assign tmp1226 = tmp1242;
    assign tmp1157 = tmp1155 ^ tmp1156;
    assign tmp1002 = tmp1018;
    assign tmp599 = tmp597 ^ tmp598;
    assign tmp1025 = {temp_15[104], temp_15[105], temp_15[106], temp_15[107], temp_15[108], temp_15[109], temp_15[110], temp_15[111]};
    assign tmp1187 = {temp_16[104], temp_16[105], temp_16[106], temp_16[107], temp_16[108], temp_16[109], temp_16[110], temp_16[111]};
    assign tmp1615 = tmp1613 ^ tmp1614;
        assign tmp421 = mem_7[tmp340];
    assign tmp957 = {temp_12[104], temp_12[105], temp_12[106], temp_12[107], temp_12[108], temp_12[109], temp_12[110], temp_12[111]};
    assign tmp1824 = {tmp1823[0], tmp1823[1], tmp1823[2], tmp1823[3], tmp1823[4], tmp1823[5], tmp1823[6], tmp1823[7]};
        assign tmp1531 = mem_7[tmp1485];
    assign tmp738 = {temp_8[16], temp_8[17], temp_8[18], temp_8[19], temp_8[20], temp_8[21], temp_8[22], temp_8[23]};
    assign b2_w7 = tmp43;
        assign tmp898 = mem_5[tmp803];
    assign tmp1335 = tmp1333 ^ tmp1334;
    assign tmp749 = {temp_9[64], temp_9[65], temp_9[66], temp_9[67], temp_9[68], temp_9[69], temp_9[70], temp_9[71]};
    assign tmp1375 = tmp1373 ^ tmp1374;
        assign tmp477 = mem_7[tmp347];
    assign tmp2244 = {tmp2243[0], tmp2243[1], tmp2243[2], tmp2243[3], tmp2243[4], tmp2243[5], tmp2243[6], tmp2243[7]};
    assign tmp1073 = tmp1071 ^ tmp1072;
    assign tmp1493 = {temp_23[40], temp_23[41], temp_23[42], temp_23[43], temp_23[44], temp_23[45], temp_23[46], temp_23[47]};
        assign tmp315 = mem_2[tmp283];
    assign tmp1654 = {temp_24[48], temp_24[49], temp_24[50], temp_24[51], temp_24[52], temp_24[53], temp_24[54], temp_24[55]};
    assign tmp1231 = tmp1247;
        assign tmp782 = mem_2[tmp750];
    assign tmp1440 = {temp_21[56], temp_21[57], temp_21[58], temp_21[59], temp_21[60], temp_21[61], temp_21[62], temp_21[63]};
    assign tmp1224 = tmp1240;
    assign tmp270 = {new_state[80], new_state[81], new_state[82], new_state[83], new_state[84], new_state[85], new_state[86], new_state[87]};
        assign tmp688 = mem_4[tmp573];
    assign temp_4 = tmp493;
    assign tmp425 = tmp423 ^ tmp424;
        assign tmp873 = mem_7[tmp799];
    assign tmp805 = {temp_11[24], temp_11[25], temp_11[26], temp_11[27], temp_11[28], temp_11[29], temp_11[30], temp_11[31]};
    assign tmp827 = tmp825 ^ tmp826;
    assign tmp1861 = tmp1859 ^ tmp1860;
    assign tmp1721 = {temp_27[56], temp_27[57], temp_27[58], temp_27[59], temp_27[60], temp_27[61], temp_27[62], temp_27[63]};
    assign tmp1605 = tmp1603 ^ tmp1604;
    assign tmp2345 = {temp_36[40], temp_36[41], temp_36[42], temp_36[43], temp_36[44], temp_36[45], temp_36[46], temp_36[47]};
    assign c1_w23 = tmp146;
    assign tmp1153 = tmp1151 ^ tmp1152;
    assign tmp2191 = tmp2228;
    assign tmp1463 = tmp1479;
        assign tmp1798 = mem_4[tmp1718];
    assign tmp530 = tmp546;
    assign tmp1105 = tmp1103 ^ tmp1104;
    assign rc4_w7 = const55_0;
    assign tmp1203 = {temp_17[112], temp_17[113], temp_17[114], temp_17[115], temp_17[116], temp_17[117], temp_17[118], temp_17[119]};
    assign tmp1799 = tmp1797 ^ tmp1798;
    assign tmp1495 = {temp_23[24], temp_23[25], temp_23[26], temp_23[27], temp_23[28], temp_23[29], temp_23[30], temp_23[31]};
    assign tmp879 = tmp877 ^ tmp878;
        assign tmp1991 = mem_7[tmp1945];
    assign tmp586 = tmp658;
    assign tmp1250 = {tmp1218, tmp1219, tmp1220, tmp1221, tmp1222, tmp1223, tmp1224, tmp1225, tmp1226, tmp1227, tmp1228, tmp1229, tmp1230, tmp1231, tmp1232, tmp1233};
    assign tmp306 = tmp322;
        assign tmp627 = mem_7[tmp567];
    assign tmp1268 = {temp_19[0], temp_19[1], temp_19[2], temp_19[3], temp_19[4], temp_19[5], temp_19[6], temp_19[7]};
    assign tmp1691 = tmp1707;
        assign tmp152 = mem_3[const151_6];
    assign tmp567 = {temp_7[88], temp_7[89], temp_7[90], temp_7[91], temp_7[92], temp_7[93], temp_7[94], temp_7[95]};
    assign tmp1272 = tmp1316;
    assign tmp1434 = {temp_21[104], temp_21[105], temp_21[106], temp_21[107], temp_21[108], temp_21[109], temp_21[110], temp_21[111]};
    assign tmp1190 = {temp_16[80], temp_16[81], temp_16[82], temp_16[83], temp_16[84], temp_16[85], temp_16[86], temp_16[87]};
    assign tmp111 = tmp110 ^ tmp86;
    assign tmp1749 = tmp1747 ^ tmp1748;
    assign tmp1597 = tmp1595 ^ tmp1596;
        assign tmp2325 = mem_7[tmp2188];
    assign tmp139 = {tmp136[8], tmp136[9], tmp136[10], tmp136[11], tmp136[12], tmp136[13], tmp136[14], tmp136[15]};
    assign tmp673 = tmp671 ^ tmp672;
        assign tmp1849 = mem_7[tmp1726];
    assign tmp2353 = {temp_37[112], temp_37[113], temp_37[114], temp_37[115], temp_37[116], temp_37[117], temp_37[118], temp_37[119]};
    assign tmp1029 = {temp_15[72], temp_15[73], temp_15[74], temp_15[75], temp_15[76], temp_15[77], temp_15[78], temp_15[79]};
    assign tmp1091 = tmp1089 ^ tmp1090;
    assign tmp964 = {temp_12[48], temp_12[49], temp_12[50], temp_12[51], temp_12[52], temp_12[53], temp_12[54], temp_12[55]};
    assign tmp476 = {tmp475[0], tmp475[1], tmp475[2], tmp475[3], tmp475[4], tmp475[5], tmp475[6], tmp475[7]};
    assign b4_w23 = tmp145;
    assign tmp1045 = tmp1110;
    assign tmp514 = {temp_5[104], temp_5[105], temp_5[106], temp_5[107], temp_5[108], temp_5[109], temp_5[110], temp_5[111]};
    assign tmp843 = tmp841 ^ tmp842;
    assign tmp751 = {temp_9[48], temp_9[49], temp_9[50], temp_9[51], temp_9[52], temp_9[53], temp_9[54], temp_9[55]};
    assign tmp87 = {tmp86[24], tmp86[25], tmp86[26], tmp86[27], tmp86[28], tmp86[29], tmp86[30], tmp86[31]};
    assign tmp1880 = {temp_28[80], temp_28[81], temp_28[82], temp_28[83], temp_28[84], temp_28[85], temp_28[86], temp_28[87]};
    assign tmp814 = tmp872;
    assign tmp1207 = {temp_17[80], temp_17[81], temp_17[82], temp_17[83], temp_17[84], temp_17[85], temp_17[86], temp_17[87]};
    assign tmp92 = {shifted_w15[24], shifted_w15[25], shifted_w15[26], shifted_w15[27], shifted_w15[28], shifted_w15[29], shifted_w15[30], shifted_w15[31]};
        assign tmp670 = mem_6[tmp574];
    assign tmp1185 = {temp_16[120], temp_16[121], temp_16[122], temp_16[123], temp_16[124], temp_16[125], temp_16[126], temp_16[127]};
        assign tmp1833 = mem_7[tmp1724];
    assign tmp1484 = {temp_23[112], temp_23[113], temp_23[114], temp_23[115], temp_23[116], temp_23[117], temp_23[118], temp_23[119]};
    assign tmp1221 = tmp1237;
    assign c2_w11 = tmp72;
    assign tmp1872 = {tmp1871[0], tmp1871[1], tmp1871[2], tmp1871[3], tmp1871[4], tmp1871[5], tmp1871[6], tmp1871[7]};
    assign tmp1633 = tmp1631 ^ tmp1632;
        assign tmp600 = mem_4[tmp566];
    assign tmp1109 = tmp1107 ^ tmp1108;
    assign tmp794 = {temp_11[112], temp_11[113], temp_11[114], temp_11[115], temp_11[116], temp_11[117], temp_11[118], temp_11[119]};
    assign tmp993 = tmp1009;
    assign tmp2231 = tmp2229 ^ tmp2230;
        assign tmp1320 = mem_6[tmp1259];
        assign tmp2330 = mem_4[tmp2187];
        assign tmp635 = mem_7[tmp568];
    assign new_5 = tmp1482;
    assign tmp2086 = {tmp2085[0], tmp2085[1], tmp2085[2], tmp2085[3], tmp2085[4], tmp2085[5], tmp2085[6], tmp2085[7]};
        assign tmp1870 = mem_4[tmp1727];
    assign tmp2368 = tmp2384;
    assign tmp575 = {temp_7[24], temp_7[25], temp_7[26], temp_7[27], temp_7[28], temp_7[29], temp_7[30], temp_7[31]};
    assign tmp1117 = tmp1115 ^ tmp1116;
    assign tmp1728 = {temp_27[0], temp_27[1], temp_27[2], temp_27[3], temp_27[4], temp_27[5], temp_27[6], temp_27[7]};
    assign tmp1102 = {tmp1101[0], tmp1101[1], tmp1101[2], tmp1101[3], tmp1101[4], tmp1101[5], tmp1101[6], tmp1101[7]};
    assign tmp393 = tmp391 ^ tmp392;
    assign tmp984 = {temp_13[24], temp_13[25], temp_13[26], temp_13[27], temp_13[28], temp_13[29], temp_13[30], temp_13[31]};
    assign tmp2321 = tmp2319 ^ tmp2320;
    assign tmp2335 = {temp_36[120], temp_36[121], temp_36[122], temp_36[123], temp_36[124], temp_36[125], temp_36[126], temp_36[127]};
    assign tmp770 = tmp786;
        assign tmp1338 = mem_4[tmp1258];
        assign tmp1566 = mem_6[tmp1487];
        assign tmp1582 = mem_6[tmp1493];
    assign tmp1585 = tmp1583 ^ tmp1584;
        assign tmp776 = mem_2[tmp744];
    assign tmp1781 = tmp1779 ^ tmp1780;
        assign tmp2290 = mem_4[tmp2182];
    assign tmp2349 = {temp_36[8], temp_36[9], temp_36[10], temp_36[11], temp_36[12], temp_36[13], temp_36[14], temp_36[15]};
    assign tmp933 = tmp931 ^ tmp932;
    assign tmp1329 = tmp1327 ^ tmp1328;
    assign tmp969 = {temp_12[8], temp_12[9], temp_12[10], temp_12[11], temp_12[12], temp_12[13], temp_12[14], temp_12[15]};
    assign tmp543 = tmp559;
    assign tmp433 = tmp431 ^ tmp432;
        assign tmp1398 = mem_5[tmp1268];
    assign concat_w19 = tmp131;
        assign tmp381 = mem_7[tmp335];
    assign tmp1348 = {tmp1347[0], tmp1347[1], tmp1347[2], tmp1347[3], tmp1347[4], tmp1347[5], tmp1347[6], tmp1347[7]};
    assign tmp978 = {temp_13[72], temp_13[73], temp_13[74], temp_13[75], temp_13[76], temp_13[77], temp_13[78], temp_13[79]};
    assign tmp2033 = tmp2031 ^ tmp2032;
    assign tmp625 = tmp623 ^ tmp624;
    assign tmp734 = {temp_8[48], temp_8[49], temp_8[50], temp_8[51], temp_8[52], temp_8[53], temp_8[54], temp_8[55]};
    assign temp_10 = tmp790;
    assign tmp1110 = {tmp1109[0], tmp1109[1], tmp1109[2], tmp1109[3], tmp1109[4], tmp1109[5], tmp1109[6], tmp1109[7]};
    assign tmp1831 = tmp1829 ^ tmp1830;
    assign tmp602 = {tmp601[0], tmp601[1], tmp601[2], tmp601[3], tmp601[4], tmp601[5], tmp601[6], tmp601[7]};
    assign tmp2360 = {temp_37[56], temp_37[57], temp_37[58], temp_37[59], temp_37[60], temp_37[61], temp_37[62], temp_37[63]};
    assign tmp244 = {shifted_w39[8], shifted_w39[9], shifted_w39[10], shifted_w39[11], shifted_w39[12], shifted_w39[13], shifted_w39[14], shifted_w39[15]};
    assign tmp303 = tmp319;
        assign tmp1777 = mem_7[tmp1717];
        assign tmp1850 = mem_5[tmp1727];
    assign b4_w27 = tmp170;
        assign tmp2293 = mem_7[tmp2184];
    assign tmp1647 = {temp_24[104], temp_24[105], temp_24[106], temp_24[107], temp_24[108], temp_24[109], temp_24[110], temp_24[111]};
    assign tmp1275 = tmp1340;
    assign tmp963 = {temp_12[56], temp_12[57], temp_12[58], temp_12[59], temp_12[60], temp_12[61], temp_12[62], temp_12[63]};
    assign tmp1219 = tmp1235;
    assign tmp2189 = tmp2212;
    assign tmp698 = {tmp697[0], tmp697[1], tmp697[2], tmp697[3], tmp697[4], tmp697[5], tmp697[6], tmp697[7]};
    assign tmp578 = {temp_7[0], temp_7[1], temp_7[2], temp_7[3], temp_7[4], temp_7[5], temp_7[6], temp_7[7]};
    assign tmp919 = tmp917 ^ tmp918;
    assign tmp655 = tmp653 ^ tmp654;
        assign tmp1328 = mem_6[tmp1260];
    assign tmp2348 = {temp_36[16], temp_36[17], temp_36[18], temp_36[19], temp_36[20], temp_36[21], temp_36[22], temp_36[23]};
    assign tmp404 = {tmp403[0], tmp403[1], tmp403[2], tmp403[3], tmp403[4], tmp403[5], tmp403[6], tmp403[7]};
        assign tmp2280 = mem_6[tmp2184];
    assign tmp2188 = {temp_35[0], temp_35[1], temp_35[2], temp_35[3], temp_35[4], temp_35[5], temp_35[6], temp_35[7]};
    assign b1_w23 = tmp142;
    assign tmp2152 = tmp2168;
    assign tmp388 = {tmp387[0], tmp387[1], tmp387[2], tmp387[3], tmp387[4], tmp387[5], tmp387[6], tmp387[7]};
    assign tmp813 = tmp864;
    assign tmp16 = {a2_w3, a3_w3, a4_w3, a1_w3};
    assign tmp296 = {temp_1[8], temp_1[9], temp_1[10], temp_1[11], temp_1[12], temp_1[13], temp_1[14], temp_1[15]};
    assign tmp1959 = tmp1982;
    assign rc1_w7 = tmp52;
    assign tmp2344 = {temp_36[48], temp_36[49], temp_36[50], temp_36[51], temp_36[52], temp_36[53], temp_36[54], temp_36[55]};
        assign tmp2082 = mem_6[tmp1958];
        assign tmp718 = mem_6[tmp576];
    assign c1_w7 = tmp46;
        assign tmp1810 = mem_5[tmp1722];
    assign tmp1594 = {tmp1593[0], tmp1593[1], tmp1593[2], tmp1593[3], tmp1593[4], tmp1593[5], tmp1593[6], tmp1593[7]};
        assign tmp908 = mem_6[tmp801];
    assign tmp11 = {aes_key[0], aes_key[1], aes_key[2], aes_key[3], aes_key[4], aes_key[5], aes_key[6], aes_key[7], aes_key[8], aes_key[9], aes_key[10], aes_key[11], aes_key[12], aes_key[13], aes_key[14], aes_key[15], aes_key[16], aes_key[17], aes_key[18], aes_key[19], aes_key[20], aes_key[21], aes_key[22], aes_key[23], aes_key[24], aes_key[25], aes_key[26], aes_key[27], aes_key[28], aes_key[29], aes_key[30], aes_key[31]};
        assign tmp2250 = mem_4[tmp2177];
    assign a3_w23 = tmp139;
    assign tmp2006 = {tmp2005[0], tmp2005[1], tmp2005[2], tmp2005[3], tmp2005[4], tmp2005[5], tmp2005[6], tmp2005[7]};
    assign tmp1689 = tmp1705;
        assign tmp1244 = mem_2[tmp1212];
        assign tmp619 = mem_7[tmp566];
    assign tmp1232 = tmp1248;
        assign tmp2302 = mem_5[tmp2186];
    assign tmp2362 = {temp_37[40], temp_37[41], temp_37[42], temp_37[43], temp_37[44], temp_37[45], temp_37[46], temp_37[47]};
    assign tmp1653 = {temp_24[56], temp_24[57], temp_24[58], temp_24[59], temp_24[60], temp_24[61], temp_24[62], temp_24[63]};
    assign c1_w39 = tmp246;
        assign tmp1249 = mem_2[tmp1217];
    assign tmp1126 = {tmp1125[0], tmp1125[1], tmp1125[2], tmp1125[3], tmp1125[4], tmp1125[5], tmp1125[6], tmp1125[7]};
        assign tmp384 = mem_6[tmp333];
    assign tmp760 = tmp776;
    assign tmp181 = {rc1_w27, rc2_w27, rc3_w27, rc4_w27};
    assign b4_w35 = tmp220;
        assign tmp2256 = mem_6[tmp2177];
    assign tmp2186 = {temp_35[16], temp_35[17], temp_35[18], temp_35[19], temp_35[20], temp_35[21], temp_35[22], temp_35[23]};
    assign tmp1851 = tmp1849 ^ tmp1850;
    assign tmp451 = tmp449 ^ tmp450;
    assign tmp1161 = tmp1159 ^ tmp1160;
        assign tmp668 = mem_5[tmp573];
    assign tmp1211 = {temp_17[48], temp_17[49], temp_17[50], temp_17[51], temp_17[52], temp_17[53], temp_17[54], temp_17[55]};
    assign temp_35 = new_2;
    assign a2_w3 = tmp13;
    assign tmp131 = {rc1_w19, rc2_w19, rc3_w19, rc4_w19};
    assign tmp2177 = {temp_35[88], temp_35[89], temp_35[90], temp_35[91], temp_35[92], temp_35[93], temp_35[94], temp_35[95]};
    assign tmp1001 = tmp1017;
    assign tmp2333 = tmp2334;
    assign tmp2340 = {temp_36[80], temp_36[81], temp_36[82], temp_36[83], temp_36[84], temp_36[85], temp_36[86], temp_36[87]};
    assign tmp1193 = {temp_16[56], temp_16[57], temp_16[58], temp_16[59], temp_16[60], temp_16[61], temp_16[62], temp_16[63]};
    assign tmp1517 = tmp1515 ^ tmp1516;
    assign tmp1735 = tmp1800;
        assign tmp1238 = mem_2[tmp1206];
    assign tmp2027 = tmp2025 ^ tmp2026;
    assign tmp43 = {shifted_w7[16], shifted_w7[17], shifted_w7[18], shifted_w7[19], shifted_w7[20], shifted_w7[21], shifted_w7[22], shifted_w7[23]};
    assign tmp298 = tmp314;
    assign tmp1760 = {tmp1759[0], tmp1759[1], tmp1759[2], tmp1759[3], tmp1759[4], tmp1759[5], tmp1759[6], tmp1759[7]};
        assign tmp2064 = mem_5[tmp1951];
    assign tmp677 = tmp675 ^ tmp676;
    assign tmp1617 = tmp1615 ^ tmp1616;
        assign tmp692 = mem_5[tmp576];
    assign tmp1483 = {temp_23[120], temp_23[121], temp_23[122], temp_23[123], temp_23[124], temp_23[125], temp_23[126], temp_23[127]};
    assign tmp212 = {tmp211[24], tmp211[25], tmp211[26], tmp211[27], tmp211[28], tmp211[29], tmp211[30], tmp211[31]};
    assign tmp1973 = tmp2094;
    assign tmp1904 = {temp_29[24], temp_29[25], temp_29[26], temp_29[27], temp_29[28], temp_29[29], temp_29[30], temp_29[31]};
    assign tmp14 = {tmp11[8], tmp11[9], tmp11[10], tmp11[11], tmp11[12], tmp11[13], tmp11[14], tmp11[15]};
    assign tmp1403 = tmp1401 ^ tmp1402;
        assign tmp2224 = mem_6[tmp2173];
    assign tmp706 = {tmp705[0], tmp705[1], tmp705[2], tmp705[3], tmp705[4], tmp705[5], tmp705[6], tmp705[7]};
    assign tmp1607 = tmp1605 ^ tmp1606;
        assign tmp598 = mem_6[tmp565];
    assign b1_w11 = tmp67;
    assign tmp83 = tmp58 ^ xor_w11;
    assign tmp125 = {c1_w19, c2_w19, c3_w19, c4_w19};
    assign tmp284 = {temp_1[104], temp_1[105], temp_1[106], temp_1[107], temp_1[108], temp_1[109], temp_1[110], temp_1[111]};
    assign tmp1763 = tmp1761 ^ tmp1762;
    assign xor_w15 = tmp107;
    assign tmp999 = tmp1015;
        assign tmp72 = mem_1[b2_w11];
    assign tmp1395 = tmp1393 ^ tmp1394;
    assign tmp981 = {temp_13[48], temp_13[49], temp_13[50], temp_13[51], temp_13[52], temp_13[53], temp_13[54], temp_13[55]};
    assign temp_37 = tmp2351;
    assign tmp1892 = {temp_29[120], temp_29[121], temp_29[122], temp_29[123], temp_29[124], temp_29[125], temp_29[126], temp_29[127]};
    assign tmp769 = tmp785;
    assign tmp2148 = tmp2164;
        assign tmp1694 = mem_2[tmp1662];
    assign tmp75 = {c1_w11, c2_w11, c3_w11, c4_w11};
    assign tmp2383 = tmp2399;
        assign tmp1635 = mem_7[tmp1498];
    assign tmp135 = tmp134 ^ tmp110;
        assign tmp2218 = mem_4[tmp2173];
        assign tmp429 = mem_7[tmp341];
        assign tmp604 = mem_5[tmp565];
    assign tmp1443 = {temp_21[32], temp_21[33], temp_21[34], temp_21[35], temp_21[36], temp_21[37], temp_21[38], temp_21[39]};
    assign tmp2173 = {temp_35[120], temp_35[121], temp_35[122], temp_35[123], temp_35[124], temp_35[125], temp_35[126], temp_35[127]};
    assign tmp592 = tmp706;
    assign tmp449 = tmp447 ^ tmp448;
    assign tmp2174 = {temp_35[112], temp_35[113], temp_35[114], temp_35[115], temp_35[116], temp_35[117], temp_35[118], temp_35[119]};
    assign tmp157 = concat_w23 ^ substituted_w23;
        assign tmp2248 = mem_6[tmp2180];
    assign tmp807 = {temp_11[8], temp_11[9], temp_11[10], temp_11[11], temp_11[12], temp_11[13], temp_11[14], temp_11[15]};
        assign tmp1168 = mem_5[tmp1038];
    assign tmp1981 = tmp1979 ^ tmp1980;
    assign tmp2110 = {temp_32[80], temp_32[81], temp_32[82], temp_32[83], temp_32[84], temp_32[85], temp_32[86], temp_32[87]};
        assign tmp1786 = mem_5[tmp1719];
    assign a4_w35 = tmp215;
        assign tmp1782 = mem_4[tmp1720];
    assign tmp848 = {tmp847[0], tmp847[1], tmp847[2], tmp847[3], tmp847[4], tmp847[5], tmp847[6], tmp847[7]};
    assign new_8 = tmp792;
        assign tmp1983 = mem_7[tmp1944];
    assign temp_14 = tmp1020;
        assign tmp1925 = mem_2[tmp1893];
    assign c4_w31 = tmp199;
        assign tmp675 = mem_7[tmp573];
        assign tmp2384 = mem_2[tmp2352];
        assign tmp454 = mem_5[tmp341];
    assign tmp2233 = tmp2231 ^ tmp2232;
    assign tmp2121 = {tmp2105, tmp2118, tmp2115, tmp2112, tmp2109, tmp2106, tmp2119, tmp2116, tmp2113, tmp2110, tmp2107, tmp2120, tmp2117, tmp2114, tmp2111, tmp2108};
    assign tmp377 = tmp375 ^ tmp376;
        assign tmp478 = mem_5[tmp348];
        assign tmp2161 = mem_2[tmp2129];
    assign tmp2364 = {temp_37[24], temp_37[25], temp_37[26], temp_37[27], temp_37[28], temp_37[29], temp_37[30], temp_37[31]};
        assign tmp1817 = mem_7[tmp1722];
    assign tmp2400 = {tmp2368, tmp2369, tmp2370, tmp2371, tmp2372, tmp2373, tmp2374, tmp2375, tmp2376, tmp2377, tmp2378, tmp2379, tmp2380, tmp2381, tmp2382, tmp2383};
        assign tmp1470 = mem_2[tmp1438];
    assign tmp1481 = {expanded_key[768], expanded_key[769], expanded_key[770], expanded_key[771], expanded_key[772], expanded_key[773], expanded_key[774], expanded_key[775], expanded_key[776], expanded_key[777], expanded_key[778], expanded_key[779], expanded_key[780], expanded_key[781], expanded_key[782], expanded_key[783], expanded_key[784], expanded_key[785], expanded_key[786], expanded_key[787], expanded_key[788], expanded_key[789], expanded_key[790], expanded_key[791], expanded_key[792], expanded_key[793], expanded_key[794], expanded_key[795], expanded_key[796], expanded_key[797], expanded_key[798], expanded_key[799], expanded_key[800], expanded_key[801], expanded_key[802], expanded_key[803], expanded_key[804], expanded_key[805], expanded_key[806], expanded_key[807], expanded_key[808], expanded_key[809], expanded_key[810], expanded_key[811], expanded_key[812], expanded_key[813], expanded_key[814], expanded_key[815], expanded_key[816], expanded_key[817], expanded_key[818], expanded_key[819], expanded_key[820], expanded_key[821], expanded_key[822], expanded_key[823], expanded_key[824], expanded_key[825], expanded_key[826], expanded_key[827], expanded_key[828], expanded_key[829], expanded_key[830], expanded_key[831], expanded_key[832], expanded_key[833], expanded_key[834], expanded_key[835], expanded_key[836], expanded_key[837], expanded_key[838], expanded_key[839], expanded_key[840], expanded_key[841], expanded_key[842], expanded_key[843], expanded_key[844], expanded_key[845], expanded_key[846], expanded_key[847], expanded_key[848], expanded_key[849], expanded_key[850], expanded_key[851], expanded_key[852], expanded_key[853], expanded_key[854], expanded_key[855], expanded_key[856], expanded_key[857], expanded_key[858], expanded_key[859], expanded_key[860], expanded_key[861], expanded_key[862], expanded_key[863], expanded_key[864], expanded_key[865], expanded_key[866], expanded_key[867], expanded_key[868], expanded_key[869], expanded_key[870], expanded_key[871], expanded_key[872], expanded_key[873], expanded_key[874], expanded_key[875], expanded_key[876], expanded_key[877], expanded_key[878], expanded_key[879], expanded_key[880], expanded_key[881], expanded_key[882], expanded_key[883], expanded_key[884], expanded_key[885], expanded_key[886], expanded_key[887], expanded_key[888], expanded_key[889], expanded_key[890], expanded_key[891], expanded_key[892], expanded_key[893], expanded_key[894], expanded_key[895]};
    assign tmp1433 = {temp_21[112], temp_21[113], temp_21[114], temp_21[115], temp_21[116], temp_21[117], temp_21[118], temp_21[119]};
    assign tmp1278 = tmp1364;
        assign tmp1374 = mem_5[tmp1261];
        assign tmp550 = mem_2[tmp518];
    assign tmp1966 = tmp2038;
        assign tmp1568 = mem_4[tmp1488];
        assign tmp672 = mem_4[tmp571];
    assign tmp200 = {c1_w31, c2_w31, c3_w31, c4_w31};
        assign tmp199 = mem_1[b4_w31];
    assign b3_w23 = tmp144;
    assign tmp2112 = {temp_32[64], temp_32[65], temp_32[66], temp_32[67], temp_32[68], temp_32[69], temp_32[70], temp_32[71]};
    assign tmp701 = tmp699 ^ tmp700;
        assign tmp1005 = mem_2[tmp973];
    assign tmp2279 = tmp2277 ^ tmp2278;
    assign tmp711 = tmp709 ^ tmp710;
    assign tmp287 = {temp_1[80], temp_1[81], temp_1[82], temp_1[83], temp_1[84], temp_1[85], temp_1[86], temp_1[87]};
    assign substituted_w31 = tmp200;
    assign tmp2089 = tmp2087 ^ tmp2088;
    assign tmp2180 = {temp_35[64], temp_35[65], temp_35[66], temp_35[67], temp_35[68], temp_35[69], temp_35[70], temp_35[71]};
    assign tmp479 = tmp477 ^ tmp478;
    assign tmp980 = {temp_13[56], temp_13[57], temp_13[58], temp_13[59], temp_13[60], temp_13[61], temp_13[62], temp_13[63]};
    assign temp_17 = tmp1201;
        assign tmp2314 = mem_4[tmp2185];
    assign tmp1513 = tmp1634;
    assign tmp40 = {tmp36[0], tmp36[1], tmp36[2], tmp36[3], tmp36[4], tmp36[5], tmp36[6], tmp36[7]};
    assign tmp979 = {temp_13[64], temp_13[65], temp_13[66], temp_13[67], temp_13[68], temp_13[69], temp_13[70], temp_13[71]};
    assign tmp1792 = {tmp1791[0], tmp1791[1], tmp1791[2], tmp1791[3], tmp1791[4], tmp1791[5], tmp1791[6], tmp1791[7]};
    assign tmp853 = tmp851 ^ tmp852;
        assign tmp551 = mem_2[tmp519];
    assign substituted_w15 = tmp100;
    assign tmp1197 = {temp_16[24], temp_16[25], temp_16[26], temp_16[27], temp_16[28], temp_16[29], temp_16[30], temp_16[31]};
    assign tmp1214 = {temp_17[24], temp_17[25], temp_17[26], temp_17[27], temp_17[28], temp_17[29], temp_17[30], temp_17[31]};
        assign tmp1590 = mem_6[tmp1494];
    assign tmp1737 = tmp1816;
    assign tmp1430 = {temp_20[0], temp_20[1], temp_20[2], temp_20[3], temp_20[4], temp_20[5], temp_20[6], temp_20[7]};
    assign tmp1897 = {temp_29[80], temp_29[81], temp_29[82], temp_29[83], temp_29[84], temp_29[85], temp_29[86], temp_29[87]};
    assign tmp965 = {temp_12[40], temp_12[41], temp_12[42], temp_12[43], temp_12[44], temp_12[45], temp_12[46], temp_12[47]};
    assign tmp114 = {tmp111[8], tmp111[9], tmp111[10], tmp111[11], tmp111[12], tmp111[13], tmp111[14], tmp111[15]};
        assign tmp608 = mem_4[tmp563];
    assign concat_w35 = tmp231;
    assign tmp1421 = {temp_20[72], temp_20[73], temp_20[74], temp_20[75], temp_20[76], temp_20[77], temp_20[78], temp_20[79]};
    assign tmp1743 = tmp1864;
    assign tmp1254 = {temp_19[112], temp_19[113], temp_19[114], temp_19[115], temp_19[116], temp_19[117], temp_19[118], temp_19[119]};
        assign tmp382 = mem_5[tmp336];
    assign tmp665 = tmp663 ^ tmp664;
        assign tmp2034 = mem_6[tmp1948];
        assign tmp432 = mem_6[tmp343];
    assign b4_w7 = tmp45;
        assign tmp2328 = mem_6[tmp2186];
    assign tmp613 = tmp611 ^ tmp612;
        assign tmp838 = mem_4[tmp793];
    assign tmp2138 = tmp2154;
    assign tmp1964 = tmp2022;
    assign tmp1291 = tmp1289 ^ tmp1290;
    assign tmp431 = tmp429 ^ tmp430;
    assign tmp2178 = {temp_35[80], temp_35[81], temp_35[82], temp_35[83], temp_35[84], temp_35[85], temp_35[86], temp_35[87]};
    assign tmp2281 = tmp2279 ^ tmp2280;
    assign tmp539 = tmp555;
        assign tmp2245 = mem_7[tmp2178];
        assign tmp96 = mem_1[b1_w15];
        assign tmp2092 = mem_4[tmp1956];
        assign tmp470 = mem_5[tmp347];
        assign tmp628 = mem_5[tmp568];
    assign tmp975 = {temp_13[96], temp_13[97], temp_13[98], temp_13[99], temp_13[100], temp_13[101], temp_13[102], temp_13[103]};
    assign tmp647 = tmp645 ^ tmp646;
        assign tmp2166 = mem_2[tmp2134];
    assign tmp591 = tmp698;
        assign tmp1286 = mem_5[tmp1254];
    assign new_state = new_11;
    assign tmp2332 = {tmp2331[0], tmp2331[1], tmp2331[2], tmp2331[3], tmp2331[4], tmp2331[5], tmp2331[6], tmp2331[7]};
    assign tmp1280 = tmp1380;
    assign tmp110 = tmp109 ^ tmp85;
    assign tmp2402 = temp_38 ^ tmp2401;
        assign tmp1858 = mem_5[tmp1728];
        assign tmp408 = mem_6[tmp340];
    assign tmp2187 = {temp_35[8], temp_35[9], temp_35[10], temp_35[11], temp_35[12], temp_35[13], temp_35[14], temp_35[15]};
    assign tmp1359 = tmp1357 ^ tmp1358;
        assign tmp1772 = mem_6[tmp1714];
        assign tmp1154 = mem_6[tmp1037];
    assign tmp2175 = {temp_35[104], temp_35[105], temp_35[106], temp_35[107], temp_35[108], temp_35[109], temp_35[110], temp_35[111]};
        assign tmp696 = mem_4[tmp578];
        assign tmp2036 = mem_4[tmp1949];
        assign tmp1532 = mem_5[tmp1486];
    assign tmp1169 = tmp1167 ^ tmp1168;
    assign tmp972 = {temp_13[120], temp_13[121], temp_13[122], temp_13[123], temp_13[124], temp_13[125], temp_13[126], temp_13[127]};
    assign tmp263 = {expanded_key[0], expanded_key[1], expanded_key[2], expanded_key[3], expanded_key[4], expanded_key[5], expanded_key[6], expanded_key[7], expanded_key[8], expanded_key[9], expanded_key[10], expanded_key[11], expanded_key[12], expanded_key[13], expanded_key[14], expanded_key[15], expanded_key[16], expanded_key[17], expanded_key[18], expanded_key[19], expanded_key[20], expanded_key[21], expanded_key[22], expanded_key[23], expanded_key[24], expanded_key[25], expanded_key[26], expanded_key[27], expanded_key[28], expanded_key[29], expanded_key[30], expanded_key[31], expanded_key[32], expanded_key[33], expanded_key[34], expanded_key[35], expanded_key[36], expanded_key[37], expanded_key[38], expanded_key[39], expanded_key[40], expanded_key[41], expanded_key[42], expanded_key[43], expanded_key[44], expanded_key[45], expanded_key[46], expanded_key[47], expanded_key[48], expanded_key[49], expanded_key[50], expanded_key[51], expanded_key[52], expanded_key[53], expanded_key[54], expanded_key[55], expanded_key[56], expanded_key[57], expanded_key[58], expanded_key[59], expanded_key[60], expanded_key[61], expanded_key[62], expanded_key[63], expanded_key[64], expanded_key[65], expanded_key[66], expanded_key[67], expanded_key[68], expanded_key[69], expanded_key[70], expanded_key[71], expanded_key[72], expanded_key[73], expanded_key[74], expanded_key[75], expanded_key[76], expanded_key[77], expanded_key[78], expanded_key[79], expanded_key[80], expanded_key[81], expanded_key[82], expanded_key[83], expanded_key[84], expanded_key[85], expanded_key[86], expanded_key[87], expanded_key[88], expanded_key[89], expanded_key[90], expanded_key[91], expanded_key[92], expanded_key[93], expanded_key[94], expanded_key[95], expanded_key[96], expanded_key[97], expanded_key[98], expanded_key[99], expanded_key[100], expanded_key[101], expanded_key[102], expanded_key[103], expanded_key[104], expanded_key[105], expanded_key[106], expanded_key[107], expanded_key[108], expanded_key[109], expanded_key[110], expanded_key[111], expanded_key[112], expanded_key[113], expanded_key[114], expanded_key[115], expanded_key[116], expanded_key[117], expanded_key[118], expanded_key[119], expanded_key[120], expanded_key[121], expanded_key[122], expanded_key[123], expanded_key[124], expanded_key[125], expanded_key[126], expanded_key[127]};
    assign tmp1391 = tmp1389 ^ tmp1390;
    assign tmp1223 = tmp1239;
        assign tmp2155 = mem_2[tmp2123];
        assign tmp2282 = mem_4[tmp2181];
        assign tmp1595 = mem_7[tmp1493];
        assign tmp1980 = mem_4[tmp1946];
        assign tmp456 = mem_6[tmp342];
        assign tmp596 = mem_5[tmp564];
    assign tmp334 = {temp_3[112], temp_3[113], temp_3[114], temp_3[115], temp_3[116], temp_3[117], temp_3[118], temp_3[119]};
    assign tmp497 = {temp_4[104], temp_4[105], temp_4[106], temp_4[107], temp_4[108], temp_4[109], temp_4[110], temp_4[111]};
    assign rc3_w39 = const254_0;
    assign tmp256 = {rc1_w39, rc2_w39, rc3_w39, rc4_w39};
    assign tmp1661 = {tmp1645, tmp1658, tmp1655, tmp1652, tmp1649, tmp1646, tmp1659, tmp1656, tmp1653, tmp1650, tmp1647, tmp1660, tmp1657, tmp1654, tmp1651, tmp1648};
        assign tmp1288 = mem_6[tmp1255];
    assign a2_w7 = tmp38;
    assign tmp1877 = {temp_28[104], temp_28[105], temp_28[106], temp_28[107], temp_28[108], temp_28[109], temp_28[110], temp_28[111]};
    assign tmp1099 = tmp1097 ^ tmp1098;
    assign tmp2276 = {tmp2275[0], tmp2275[1], tmp2275[2], tmp2275[3], tmp2275[4], tmp2275[5], tmp2275[6], tmp2275[7]};
    assign tmp395 = tmp393 ^ tmp394;
        assign tmp1518 = mem_6[tmp1485];
        assign tmp1060 = mem_4[tmp1026];
        assign tmp1006 = mem_2[tmp974];
    assign tmp1033 = {temp_15[40], temp_15[41], temp_15[42], temp_15[43], temp_15[44], temp_15[45], temp_15[46], temp_15[47]};
    assign tmp1177 = tmp1175 ^ tmp1176;
    assign tmp1425 = {temp_20[40], temp_20[41], temp_20[42], temp_20[43], temp_20[44], temp_20[45], temp_20[46], temp_20[47]};
    assign tmp536 = tmp552;
        assign tmp1611 = mem_7[tmp1495];
    assign tmp66 = {a2_w11, a3_w11, a4_w11, a1_w11};
    assign tmp531 = tmp547;
    assign tmp525 = {temp_5[16], temp_5[17], temp_5[18], temp_5[19], temp_5[20], temp_5[21], temp_5[22], temp_5[23]};
        assign tmp2213 = mem_7[tmp2174];
    assign tmp2057 = tmp2055 ^ tmp2056;
    assign c3_w39 = tmp248;
    assign tmp1651 = {temp_24[72], temp_24[73], temp_24[74], temp_24[75], temp_24[76], temp_24[77], temp_24[78], temp_24[79]};
    assign tmp855 = tmp853 ^ tmp854;
        assign tmp881 = mem_7[tmp800];
    assign tmp2106 = {temp_32[112], temp_32[113], temp_32[114], temp_32[115], temp_32[116], temp_32[117], temp_32[118], temp_32[119]};
    assign b3_w7 = tmp44;
    assign tmp2376 = tmp2392;
    assign shifted_w7 = tmp41;
    assign tmp1800 = {tmp1799[0], tmp1799[1], tmp1799[2], tmp1799[3], tmp1799[4], tmp1799[5], tmp1799[6], tmp1799[7]};
    assign tmp1042 = tmp1086;
        assign tmp392 = mem_6[tmp334];
        assign tmp2399 = mem_2[tmp2367];
    assign tmp2212 = {tmp2211[0], tmp2211[1], tmp2211[2], tmp2211[3], tmp2211[4], tmp2211[5], tmp2211[6], tmp2211[7]};
    assign tmp1508 = tmp1594;
        assign tmp1695 = mem_2[tmp1663];
    assign tmp974 = {temp_13[104], temp_13[105], temp_13[106], temp_13[107], temp_13[108], temp_13[109], temp_13[110], temp_13[111]};
    assign tmp997 = tmp1013;
    assign tmp1787 = tmp1785 ^ tmp1786;
    assign shifted_w11 = tmp66;
        assign tmp707 = mem_7[tmp577];
    assign tmp299 = tmp315;
    assign new_9 = tmp562;
    assign tmp991 = tmp1007;
    assign tmp2136 = {temp_33[8], temp_33[9], temp_33[10], temp_33[11], temp_33[12], temp_33[13], temp_33[14], temp_33[15]};
    assign tmp1673 = {temp_25[32], temp_25[33], temp_25[34], temp_25[35], temp_25[36], temp_25[37], temp_25[38], temp_25[39]};
    assign tmp1726 = {temp_27[16], temp_27[17], temp_27[18], temp_27[19], temp_27[20], temp_27[21], temp_27[22], temp_27[23]};
    assign tmp2022 = {tmp2021[0], tmp2021[1], tmp2021[2], tmp2021[3], tmp2021[4], tmp2021[5], tmp2021[6], tmp2021[7]};
    assign tmp1171 = tmp1169 ^ tmp1170;
    assign tmp1808 = {tmp1807[0], tmp1807[1], tmp1807[2], tmp1807[3], tmp1807[4], tmp1807[5], tmp1807[6], tmp1807[7]};
    assign tmp1300 = {tmp1299[0], tmp1299[1], tmp1299[2], tmp1299[3], tmp1299[4], tmp1299[5], tmp1299[6], tmp1299[7]};
    assign tmp371 = tmp369 ^ tmp370;
    assign tmp621 = tmp619 ^ tmp620;
    assign tmp2101 = tmp2099 ^ tmp2100;
        assign tmp378 = mem_4[tmp333];
    assign tmp1077 = tmp1075 ^ tmp1076;
    assign tmp118 = {shifted_w19[16], shifted_w19[17], shifted_w19[18], shifted_w19[19], shifted_w19[20], shifted_w19[21], shifted_w19[22], shifted_w19[23]};
    assign tmp2329 = tmp2327 ^ tmp2328;
        assign tmp434 = mem_4[tmp344];
    assign tmp156 = {rc1_w23, rc2_w23, rc3_w23, rc4_w23};
    assign tmp187 = {tmp186[24], tmp186[25], tmp186[26], tmp186[27], tmp186[28], tmp186[29], tmp186[30], tmp186[31]};
        assign tmp469 = mem_7[tmp346];
    assign tmp391 = tmp389 ^ tmp390;
    assign tmp601 = tmp599 ^ tmp600;
    assign tmp1388 = {tmp1387[0], tmp1387[1], tmp1387[2], tmp1387[3], tmp1387[4], tmp1387[5], tmp1387[6], tmp1387[7]};
    assign tmp1883 = {temp_28[56], temp_28[57], temp_28[58], temp_28[59], temp_28[60], temp_28[61], temp_28[62], temp_28[63]};
        assign tmp1704 = mem_2[tmp1672];
    assign b3_w3 = tmp19;
    assign tmp529 = tmp545;
    assign tmp504 = {temp_4[48], temp_4[49], temp_4[50], temp_4[51], temp_4[52], temp_4[53], temp_4[54], temp_4[55]};
    assign tmp1791 = tmp1789 ^ tmp1790;
        assign tmp1055 = mem_7[tmp1023];
    assign tmp348 = {temp_3[0], temp_3[1], temp_3[2], temp_3[3], temp_3[4], temp_3[5], temp_3[6], temp_3[7]};
    assign tmp349 = tmp372;
    assign tmp300 = tmp316;
        assign tmp1140 = mem_4[tmp1032];
    assign tmp1252 = temp_18 ^ tmp1251;
        assign tmp544 = mem_2[tmp512];
    assign tmp1217 = {temp_17[0], temp_17[1], temp_17[2], temp_17[3], temp_17[4], temp_17[5], temp_17[6], temp_17[7]};
        assign tmp2398 = mem_2[tmp2366];
    assign tmp542 = tmp558;
    assign tmp1445 = {temp_21[16], temp_21[17], temp_21[18], temp_21[19], temp_21[20], temp_21[21], temp_21[22], temp_21[23]};
        assign tmp2286 = mem_5[tmp2184];
    assign tmp1367 = tmp1365 ^ tmp1366;
        assign tmp616 = mem_4[tmp564];
    assign tmp1316 = {tmp1315[0], tmp1315[1], tmp1315[2], tmp1315[3], tmp1315[4], tmp1315[5], tmp1315[6], tmp1315[7]};
    assign a4_w7 = tmp40;
        assign tmp1834 = mem_5[tmp1721];
    assign tmp523 = {temp_5[32], temp_5[33], temp_5[34], temp_5[35], temp_5[36], temp_5[37], temp_5[38], temp_5[39]};
        assign tmp1116 = mem_4[tmp1029];
    assign tmp573 = {temp_7[40], temp_7[41], temp_7[42], temp_7[43], temp_7[44], temp_7[45], temp_7[46], temp_7[47]};
    assign tmp159 = tmp158 ^ tmp134;
    assign tmp1461 = tmp1477;
    assign tmp2331 = tmp2329 ^ tmp2330;
        assign tmp1700 = mem_2[tmp1668];
        assign tmp664 = mem_4[tmp574];
        assign tmp1015 = mem_2[tmp983];
    assign rc1_w19 = tmp127;
    assign temp_28 = tmp1873;
        assign tmp894 = mem_4[tmp804];
    assign tmp499 = {temp_4[88], temp_4[89], temp_4[90], temp_4[91], temp_4[92], temp_4[93], temp_4[94], temp_4[95]};
    assign tmp723 = tmp724;
    assign tmp1199 = {temp_16[8], temp_16[9], temp_16[10], temp_16[11], temp_16[12], temp_16[13], temp_16[14], temp_16[15]};
    assign tmp444 = {tmp443[0], tmp443[1], tmp443[2], tmp443[3], tmp443[4], tmp443[5], tmp443[6], tmp443[7]};
    assign tmp182 = concat_w27 ^ substituted_w27;
    assign tmp2075 = tmp2073 ^ tmp2074;
    assign tmp484 = {tmp483[0], tmp483[1], tmp483[2], tmp483[3], tmp483[4], tmp483[5], tmp483[6], tmp483[7]};
    assign tmp290 = {temp_1[56], temp_1[57], temp_1[58], temp_1[59], temp_1[60], temp_1[61], temp_1[62], temp_1[63]};
    assign tmp259 = tmp258 ^ tmp234;
        assign tmp1809 = mem_7[tmp1721];
        assign tmp2157 = mem_2[tmp2125];
        assign tmp1598 = mem_6[tmp1491];
        assign tmp2087 = mem_7[tmp1957];
    assign tmp1453 = tmp1469;
    assign tmp1837 = tmp1835 ^ tmp1836;
    assign tmp501 = {temp_4[72], temp_4[73], temp_4[74], temp_4[75], temp_4[76], temp_4[77], temp_4[78], temp_4[79]};
        assign tmp910 = mem_4[tmp802];
        assign tmp1381 = mem_7[tmp1265];
    assign tmp281 = {tmp265, tmp278, tmp275, tmp272, tmp269, tmp266, tmp279, tmp276, tmp273, tmp270, tmp267, tmp280, tmp277, tmp274, tmp271, tmp268};
        assign tmp318 = mem_2[tmp286];
    assign a1_w3 = tmp12;
    assign tmp1218 = tmp1234;
    assign tmp1989 = tmp1987 ^ tmp1988;
    assign tmp1504 = tmp1562;
        assign tmp849 = mem_7[tmp796];
        assign tmp1624 = mem_4[tmp1495];
        assign tmp710 = mem_6[tmp575];
    assign tmp568 = {temp_7[80], temp_7[81], temp_7[82], temp_7[83], temp_7[84], temp_7[85], temp_7[86], temp_7[87]};
        assign tmp2285 = mem_7[tmp2183];
        assign tmp222 = mem_1[b2_w35];
    assign tmp1050 = tmp1150;
    assign c3_w15 = tmp98;
        assign tmp1302 = mem_5[tmp1256];
    assign tmp1271 = tmp1308;
        assign tmp2060 = mem_4[tmp1952];
        assign tmp1466 = mem_2[tmp1434];
        assign tmp406 = mem_5[tmp339];
        assign tmp651 = mem_7[tmp570];
        assign tmp950 = mem_4[tmp807];
    assign tmp2260 = {tmp2259[0], tmp2259[1], tmp2259[2], tmp2259[3], tmp2259[4], tmp2259[5], tmp2259[6], tmp2259[7]};
    assign tmp823 = tmp944;
    assign tmp1759 = tmp1757 ^ tmp1758;
    assign temp_9 = tmp741;
    assign tmp804 = {temp_11[32], temp_11[33], temp_11[34], temp_11[35], temp_11[36], temp_11[37], temp_11[38], temp_11[39]};
    assign tmp1500 = tmp1530;
    assign tmp732 = {temp_8[64], temp_8[65], temp_8[66], temp_8[67], temp_8[68], temp_8[69], temp_8[70], temp_8[71]};
    assign tmp893 = tmp891 ^ tmp892;
    assign tmp1670 = {temp_25[56], temp_25[57], temp_25[58], temp_25[59], temp_25[60], temp_25[61], temp_25[62], temp_25[63]};
    assign a2_w39 = tmp238;
        assign tmp1464 = mem_2[tmp1432];
    assign tmp1257 = {temp_19[88], temp_19[89], temp_19[90], temp_19[91], temp_19[92], temp_19[93], temp_19[94], temp_19[95]};
        assign tmp1584 = mem_4[tmp1494];
        assign tmp686 = mem_6[tmp572];
    assign new_7 = tmp1022;
        assign tmp1706 = mem_2[tmp1674];
        assign tmp870 = mem_4[tmp797];
    assign tmp1908 = tmp1924;
    assign tmp973 = {temp_13[112], temp_13[113], temp_13[114], temp_13[115], temp_13[116], temp_13[117], temp_13[118], temp_13[119]};
    assign temp_1 = tmp281;
        assign tmp2088 = mem_5[tmp1958];
    assign tmp20 = {shifted_w3[0], shifted_w3[1], shifted_w3[2], shifted_w3[3], shifted_w3[4], shifted_w3[5], shifted_w3[6], shifted_w3[7]};
    assign xor_w31 = tmp207;
        assign tmp482 = mem_4[tmp346];
        assign tmp702 = mem_6[tmp578];
        assign tmp2080 = mem_5[tmp1957];
    assign tmp1567 = tmp1565 ^ tmp1566;
        assign tmp1476 = mem_2[tmp1444];
    assign tmp1902 = {temp_29[40], temp_29[41], temp_29[42], temp_29[43], temp_29[44], temp_29[45], temp_29[46], temp_29[47]};
    assign tmp1577 = tmp1575 ^ tmp1576;
        assign tmp430 = mem_5[tmp342];
    assign tmp1684 = tmp1700;
    assign b1_w27 = tmp167;
    assign tmp2147 = tmp2163;
    assign tmp307 = tmp323;
    assign tmp2219 = tmp2217 ^ tmp2218;
    assign tmp1075 = tmp1073 ^ tmp1074;
    assign tmp1401 = tmp1399 ^ tmp1400;
    assign tmp1819 = tmp1817 ^ tmp1818;
        assign tmp1548 = mem_5[tmp1488];
    assign tmp1879 = {temp_28[88], temp_28[89], temp_28[90], temp_28[91], temp_28[92], temp_28[93], temp_28[94], temp_28[95]};
    assign tmp824 = tmp952;
    assign tmp800 = {temp_11[64], temp_11[65], temp_11[66], temp_11[67], temp_11[68], temp_11[69], temp_11[70], temp_11[71]};
    assign tmp1910 = tmp1926;
        assign tmp2040 = mem_5[tmp1952];
    assign tmp821 = tmp928;
        assign tmp700 = mem_5[tmp577];
    assign tmp837 = tmp835 ^ tmp836;
    assign tmp1387 = tmp1385 ^ tmp1386;
        assign tmp376 = mem_6[tmp336];
    assign tmp1768 = {tmp1767[0], tmp1767[1], tmp1767[2], tmp1767[3], tmp1767[4], tmp1767[5], tmp1767[6], tmp1767[7]};
    assign tmp61 = tmp60 ^ tmp36;
        assign tmp1138 = mem_6[tmp1031];
    assign c4_w39 = tmp249;
    assign tmp2179 = {temp_35[72], temp_35[73], temp_35[74], temp_35[75], temp_35[76], temp_35[77], temp_35[78], temp_35[79]};
    assign tmp1123 = tmp1121 ^ tmp1122;
        assign tmp2162 = mem_2[tmp2130];
        assign tmp1172 = mem_4[tmp1036];
    assign tmp258 = tmp233 ^ xor_w39;
    assign tmp225 = {c1_w35, c2_w35, c3_w35, c4_w35};
    assign tmp2341 = {temp_36[72], temp_36[73], temp_36[74], temp_36[75], temp_36[76], temp_36[77], temp_36[78], temp_36[79]};
    assign tmp1641 = tmp1639 ^ tmp1640;
        assign tmp1474 = mem_2[tmp1442];
    assign tmp143 = {shifted_w23[16], shifted_w23[17], shifted_w23[18], shifted_w23[19], shifted_w23[20], shifted_w23[21], shifted_w23[22], shifted_w23[23]};
    assign tmp184 = tmp183 ^ tmp159;
    assign tmp2025 = tmp2023 ^ tmp2024;
    assign tmp2107 = {temp_32[104], temp_32[105], temp_32[106], temp_32[107], temp_32[108], temp_32[109], temp_32[110], temp_32[111]};
        assign tmp1933 = mem_2[tmp1901];
    assign tmp757 = {temp_9[0], temp_9[1], temp_9[2], temp_9[3], temp_9[4], temp_9[5], temp_9[6], temp_9[7]};
    assign tmp1047 = tmp1126;
    assign concat_w31 = tmp206;
        assign tmp1812 = mem_6[tmp1723];
    assign rc2_w39 = const253_0;
    assign tmp756 = {temp_9[8], temp_9[9], temp_9[10], temp_9[11], temp_9[12], temp_9[13], temp_9[14], temp_9[15]};
    assign a2_w11 = tmp63;
    assign tmp983 = {temp_13[32], temp_13[33], temp_13[34], temp_13[35], temp_13[36], temp_13[37], temp_13[38], temp_13[39]};
    assign tmp1258 = {temp_19[80], temp_19[81], temp_19[82], temp_19[83], temp_19[84], temp_19[85], temp_19[86], temp_19[87]};
    assign tmp2185 = {temp_35[24], temp_35[25], temp_35[26], temp_35[27], temp_35[28], temp_35[29], temp_35[30], temp_35[31]};
    assign tmp1970 = tmp2070;
        assign tmp2269 = mem_7[tmp2181];
    assign tmp1602 = {tmp1601[0], tmp1601[1], tmp1601[2], tmp1601[3], tmp1601[4], tmp1601[5], tmp1601[6], tmp1601[7]};
    assign tmp1795 = tmp1793 ^ tmp1794;
    assign tmp492 = {tmp491[0], tmp491[1], tmp491[2], tmp491[3], tmp491[4], tmp491[5], tmp491[6], tmp491[7]};
    assign tmp761 = tmp777;
    assign tmp1715 = {temp_27[104], temp_27[105], temp_27[106], temp_27[107], temp_27[108], temp_27[109], temp_27[110], temp_27[111]};
    assign tmp236 = tmp235 ^ tmp211;
    assign b4_w15 = tmp95;
        assign tmp1400 = mem_6[tmp1265];
    assign tmp515 = {temp_5[96], temp_5[97], temp_5[98], temp_5[99], temp_5[100], temp_5[101], temp_5[102], temp_5[103]};
    assign tmp457 = tmp455 ^ tmp456;
        assign tmp2254 = mem_5[tmp2180];
    assign tmp158 = tmp133 ^ xor_w23;
    assign tmp1951 = {temp_31[56], temp_31[57], temp_31[58], temp_31[59], temp_31[60], temp_31[61], temp_31[62], temp_31[63]};
    assign tmp2295 = tmp2293 ^ tmp2294;
    assign tmp107 = concat_w15 ^ substituted_w15;
    assign tmp790 = {tmp758, tmp759, tmp760, tmp761, tmp762, tmp763, tmp764, tmp765, tmp766, tmp767, tmp768, tmp769, tmp770, tmp771, tmp772, tmp773};
    assign tmp755 = {temp_9[16], temp_9[17], temp_9[18], temp_9[19], temp_9[20], temp_9[21], temp_9[22], temp_9[23]};
    assign tmp2146 = tmp2162;
    assign tmp1676 = {temp_25[8], temp_25[9], temp_25[10], temp_25[11], temp_25[12], temp_25[13], temp_25[14], temp_25[15]};
    assign tmp1771 = tmp1769 ^ tmp1770;
    assign tmp1783 = tmp1781 ^ tmp1782;
    assign tmp1455 = tmp1471;
        assign tmp865 = mem_7[tmp798];
        assign tmp547 = mem_2[tmp515];
    assign temp_13 = tmp971;
        assign tmp1558 = mem_6[tmp1490];
    assign a1_w15 = tmp87;
    assign tmp1439 = {temp_21[64], temp_21[65], temp_21[66], temp_21[67], temp_21[68], temp_21[69], temp_21[70], temp_21[71]};
        assign tmp854 = mem_4[tmp795];
    assign tmp912 = {tmp911[0], tmp911[1], tmp911[2], tmp911[3], tmp911[4], tmp911[5], tmp911[6], tmp911[7]};
    assign tmp511 = {tmp495, tmp508, tmp505, tmp502, tmp499, tmp496, tmp509, tmp506, tmp503, tmp500, tmp497, tmp510, tmp507, tmp504, tmp501, tmp498};
    assign tmp279 = {new_state[8], new_state[9], new_state[10], new_state[11], new_state[12], new_state[13], new_state[14], new_state[15]};
    assign tmp1052 = tmp1166;
    assign tmp1739 = tmp1832;
    assign tmp1451 = tmp1467;
    assign tmp1107 = tmp1105 ^ tmp1106;
    assign tmp2059 = tmp2057 ^ tmp2058;
    assign tmp379 = tmp377 ^ tmp378;
    assign tmp1955 = {temp_31[24], temp_31[25], temp_31[26], temp_31[27], temp_31[28], temp_31[29], temp_31[30], temp_31[31]};
    assign tmp1442 = {temp_21[40], temp_21[41], temp_21[42], temp_21[43], temp_21[44], temp_21[45], temp_21[46], temp_21[47]};
    assign a1_w7 = tmp37;
        assign tmp652 = mem_5[tmp567];
    assign tmp2211 = tmp2209 ^ tmp2210;
        assign tmp1152 = mem_5[tmp1036];
    assign tmp2292 = {tmp2291[0], tmp2291[1], tmp2291[2], tmp2291[3], tmp2291[4], tmp2291[5], tmp2291[6], tmp2291[7]};
    assign tmp1565 = tmp1563 ^ tmp1564;
    assign tmp1886 = {temp_28[32], temp_28[33], temp_28[34], temp_28[35], temp_28[36], temp_28[37], temp_28[38], temp_28[39]};
    assign tmp1133 = tmp1131 ^ tmp1132;
        assign tmp683 = mem_7[tmp574];
        assign tmp438 = mem_5[tmp343];
    assign tmp956 = {temp_12[112], temp_12[113], temp_12[114], temp_12[115], temp_12[116], temp_12[117], temp_12[118], temp_12[119]};
    assign tmp566 = {temp_7[96], temp_7[97], temp_7[98], temp_7[99], temp_7[100], temp_7[101], temp_7[102], temp_7[103]};
    assign rc4_w3 = const30_0;
    assign tmp1385 = tmp1383 ^ tmp1384;
        assign tmp556 = mem_2[tmp524];
    assign tmp1459 = tmp1475;
        assign tmp900 = mem_6[tmp804];
    assign tmp1686 = tmp1702;
    assign tmp565 = {temp_7[104], temp_7[105], temp_7[106], temp_7[107], temp_7[108], temp_7[109], temp_7[110], temp_7[111]};
        assign tmp1860 = mem_6[tmp1725];
    assign tmp1888 = {temp_28[16], temp_28[17], temp_28[18], temp_28[19], temp_28[20], temp_28[21], temp_28[22], temp_28[23]};
    assign tmp1960 = tmp1990;
    assign temp_36 = tmp2333;
    assign tmp650 = {tmp649[0], tmp649[1], tmp649[2], tmp649[3], tmp649[4], tmp649[5], tmp649[6], tmp649[7]};
        assign tmp549 = mem_2[tmp517];
        assign tmp886 = mem_4[tmp799];
    assign tmp1494 = {temp_23[32], temp_23[33], temp_23[34], temp_23[35], temp_23[36], temp_23[37], temp_23[38], temp_23[39]};
    assign tmp812 = tmp856;
    assign tmp88 = {tmp86[16], tmp86[17], tmp86[18], tmp86[19], tmp86[20], tmp86[21], tmp86[22], tmp86[23]};
    assign tmp359 = tmp452;
    assign tmp1537 = tmp1535 ^ tmp1536;
    assign tmp206 = {rc1_w31, rc2_w31, rc3_w31, rc4_w31};
    assign tmp185 = tmp184 ^ tmp160;
        assign tmp558 = mem_2[tmp526];
    assign c1_w31 = tmp196;
        assign tmp1935 = mem_2[tmp1903];
        assign tmp1468 = mem_2[tmp1436];
    assign tmp1174 = {tmp1173[0], tmp1173[1], tmp1173[2], tmp1173[3], tmp1173[4], tmp1173[5], tmp1173[6], tmp1173[7]};
        assign tmp1560 = mem_4[tmp1487];
        assign tmp1555 = mem_7[tmp1488];
        assign tmp71 = mem_1[b1_w11];
    assign tmp240 = {tmp236[0], tmp236[1], tmp236[2], tmp236[3], tmp236[4], tmp236[5], tmp236[6], tmp236[7]};
    assign tmp163 = {tmp161[16], tmp161[17], tmp161[18], tmp161[19], tmp161[20], tmp161[21], tmp161[22], tmp161[23]};
    assign tmp1273 = tmp1324;
        assign tmp1804 = mem_6[tmp1718];
        assign tmp319 = mem_2[tmp287];
    assign tmp39 = {tmp36[8], tmp36[9], tmp36[10], tmp36[11], tmp36[12], tmp36[13], tmp36[14], tmp36[15]};
    assign tmp2061 = tmp2059 ^ tmp2060;
    assign tmp2380 = tmp2396;
    assign tmp709 = tmp707 ^ tmp708;
        assign tmp1120 = mem_5[tmp1032];
    assign tmp1519 = tmp1517 ^ tmp1518;
    assign tmp1024 = {temp_15[112], temp_15[113], temp_15[114], temp_15[115], temp_15[116], temp_15[117], temp_15[118], temp_15[119]};
    assign tmp312 = tmp328;
    assign tmp1538 = {tmp1537[0], tmp1537[1], tmp1537[2], tmp1537[3], tmp1537[4], tmp1537[5], tmp1537[6], tmp1537[7]};
    assign tmp487 = tmp485 ^ tmp486;
    assign tmp1642 = {tmp1641[0], tmp1641[1], tmp1641[2], tmp1641[3], tmp1641[4], tmp1641[5], tmp1641[6], tmp1641[7]};
    assign tmp2370 = tmp2386;
    assign tmp911 = tmp909 ^ tmp910;
        assign tmp413 = mem_7[tmp339];
    assign rc3_w19 = const129_0;
    assign tmp1655 = {temp_24[40], temp_24[41], temp_24[42], temp_24[43], temp_24[44], temp_24[45], temp_24[46], temp_24[47]};
    assign tmp1284 = tmp1412;
        assign tmp937 = mem_7[tmp807];
        assign tmp488 = mem_6[tmp346];
    assign tmp1480 = {tmp1448, tmp1449, tmp1450, tmp1451, tmp1452, tmp1453, tmp1454, tmp1455, tmp1456, tmp1457, tmp1458, tmp1459, tmp1460, tmp1461, tmp1462, tmp1463};
    assign tmp1971 = tmp2078;
    assign tmp2355 = {temp_37[96], temp_37[97], temp_37[98], temp_37[99], temp_37[100], temp_37[101], temp_37[102], temp_37[103]};
        assign tmp2242 = mem_4[tmp2180];
        assign tmp365 = mem_7[tmp333];
        assign tmp922 = mem_5[tmp806];
    assign rc1_w27 = tmp177;
    assign tmp798 = {temp_11[80], temp_11[81], temp_11[82], temp_11[83], temp_11[84], temp_11[85], temp_11[86], temp_11[87]};
    assign tmp241 = {a2_w39, a3_w39, a4_w39, a1_w39};
        assign tmp1294 = mem_5[tmp1255];
    assign b4_w39 = tmp245;
    assign tmp351 = tmp388;
    assign tmp67 = {shifted_w11[24], shifted_w11[25], shifted_w11[26], shifted_w11[27], shifted_w11[28], shifted_w11[29], shifted_w11[30], shifted_w11[31]};
    assign tmp1660 = {temp_24[0], temp_24[1], temp_24[2], temp_24[3], temp_24[4], temp_24[5], temp_24[6], temp_24[7]};
    assign tmp481 = tmp479 ^ tmp480;
    assign c4_w23 = tmp149;
        assign tmp846 = mem_4[tmp794];
        assign tmp834 = mem_5[tmp795];
    assign tmp1502 = tmp1546;
    assign tmp427 = tmp425 ^ tmp426;
    assign tmp1954 = {temp_31[32], temp_31[33], temp_31[34], temp_31[35], temp_31[36], temp_31[37], temp_31[38], temp_31[39]};
    assign tmp1855 = tmp1853 ^ tmp1854;
        assign tmp1469 = mem_2[tmp1437];
    assign tmp954 = {tmp809, tmp810, tmp811, tmp812, tmp813, tmp814, tmp815, tmp816, tmp817, tmp818, tmp819, tmp820, tmp821, tmp822, tmp823, tmp824};
    assign tmp887 = tmp885 ^ tmp886;
        assign tmp1366 = mem_5[tmp1264];
    assign tmp339 = {temp_3[72], temp_3[73], temp_3[74], temp_3[75], temp_3[76], temp_3[77], temp_3[78], temp_3[79]};
        assign tmp2272 = mem_6[tmp2183];
    assign tmp1202 = {temp_17[120], temp_17[121], temp_17[122], temp_17[123], temp_17[124], temp_17[125], temp_17[126], temp_17[127]};
    assign tmp909 = tmp907 ^ tmp908;
        assign tmp1758 = mem_4[tmp1713];
    assign tmp1446 = {temp_21[8], temp_21[9], temp_21[10], temp_21[11], temp_21[12], temp_21[13], temp_21[14], temp_21[15]};
    assign a2_w23 = tmp138;
        assign tmp691 = mem_7[tmp575];
    assign tmp1345 = tmp1343 ^ tmp1344;
    assign c2_w31 = tmp197;
    assign tmp532 = tmp548;
        assign tmp1988 = mem_4[tmp1943];
        assign tmp1619 = mem_7[tmp1496];
        assign tmp1926 = mem_2[tmp1894];
        assign tmp787 = mem_2[tmp755];
    assign tmp1255 = {temp_19[104], temp_19[105], temp_19[106], temp_19[107], temp_19[108], temp_19[109], temp_19[110], temp_19[111]};
    assign tmp1535 = tmp1533 ^ tmp1534;
    assign tmp2142 = tmp2158;
    assign tmp1887 = {temp_28[24], temp_28[25], temp_28[26], temp_28[27], temp_28[28], temp_28[29], temp_28[30], temp_28[31]};
    assign temp_16 = tmp1183;
    assign tmp742 = {temp_9[120], temp_9[121], temp_9[122], temp_9[123], temp_9[124], temp_9[125], temp_9[126], temp_9[127]};
    assign tmp1189 = {temp_16[88], temp_16[89], temp_16[90], temp_16[91], temp_16[92], temp_16[93], temp_16[94], temp_16[95]};
    assign tmp1195 = {temp_16[40], temp_16[41], temp_16[42], temp_16[43], temp_16[44], temp_16[45], temp_16[46], temp_16[47]};
        assign tmp1814 = mem_4[tmp1724];
    assign tmp1028 = {temp_15[80], temp_15[81], temp_15[82], temp_15[83], temp_15[84], temp_15[85], temp_15[86], temp_15[87]};
    assign tmp1525 = tmp1523 ^ tmp1524;
    assign temp_8 = tmp723;
        assign tmp906 = mem_5[tmp804];
    assign tmp1593 = tmp1591 ^ tmp1592;
    assign tmp217 = {shifted_w35[24], shifted_w35[25], shifted_w35[26], shifted_w35[27], shifted_w35[28], shifted_w35[29], shifted_w35[30], shifted_w35[31]};
    assign a3_w3 = tmp14;
        assign tmp1934 = mem_2[tmp1902];
        assign tmp2296 = mem_6[tmp2182];
    assign b1_w3 = tmp17;
    assign c2_w27 = tmp172;
    assign tmp1431 = {tmp1415, tmp1428, tmp1425, tmp1422, tmp1419, tmp1416, tmp1429, tmp1426, tmp1423, tmp1420, tmp1417, tmp1430, tmp1427, tmp1424, tmp1421, tmp1418};
    assign tmp883 = tmp881 ^ tmp882;
        assign tmp1547 = mem_7[tmp1487];
        assign tmp171 = mem_1[b1_w27];
        assign tmp918 = mem_4[tmp803];
    assign tmp952 = {tmp951[0], tmp951[1], tmp951[2], tmp951[3], tmp951[4], tmp951[5], tmp951[6], tmp951[7]};
    assign temp_7 = new_9;
    assign tmp989 = tmp1005;
    assign tmp1230 = tmp1246;
    assign tmp1196 = {temp_16[32], temp_16[33], temp_16[34], temp_16[35], temp_16[36], temp_16[37], temp_16[38], temp_16[39]};
    assign tmp1097 = tmp1095 ^ tmp1096;
    assign tmp721 = tmp719 ^ tmp720;
    assign tmp816 = tmp888;
        assign tmp1526 = mem_6[tmp1486];
    assign tmp537 = tmp553;
    assign tmp1779 = tmp1777 ^ tmp1778;
    assign tmp141 = {a2_w23, a3_w23, a4_w23, a1_w23};
    assign tmp815 = tmp880;
    assign tmp356 = tmp428;
        assign tmp1596 = mem_5[tmp1494];
    assign tmp1496 = {temp_23[16], temp_23[17], temp_23[18], temp_23[19], temp_23[20], temp_23[21], temp_23[22], temp_23[23]};
        assign tmp1076 = mem_4[tmp1024];
        assign tmp1012 = mem_2[tmp980];
    assign tmp1885 = {temp_28[40], temp_28[41], temp_28[42], temp_28[43], temp_28[44], temp_28[45], temp_28[46], temp_28[47]};
    assign tmp1634 = {tmp1633[0], tmp1633[1], tmp1633[2], tmp1633[3], tmp1633[4], tmp1633[5], tmp1633[6], tmp1633[7]};
        assign tmp394 = mem_4[tmp335];
    assign a4_w11 = tmp65;
        assign tmp2312 = mem_6[tmp2188];
    assign tmp1418 = {temp_20[96], temp_20[97], temp_20[98], temp_20[99], temp_20[100], temp_20[101], temp_20[102], temp_20[103]};
    assign tmp1462 = tmp1478;
    assign tmp64 = {tmp61[8], tmp61[9], tmp61[10], tmp61[11], tmp61[12], tmp61[13], tmp61[14], tmp61[15]};
    assign tmp1420 = {temp_20[80], temp_20[81], temp_20[82], temp_20[83], temp_20[84], temp_20[85], temp_20[86], temp_20[87]};
    assign tmp689 = tmp687 ^ tmp688;
    assign tmp538 = tmp554;
        assign tmp196 = mem_1[b1_w31];
        assign tmp1290 = mem_4[tmp1256];
        assign tmp929 = mem_7[tmp806];
        assign tmp2393 = mem_2[tmp2361];
    assign tmp1688 = tmp1704;
        assign tmp1638 = mem_6[tmp1496];
    assign tmp1733 = tmp1784;
        assign tmp546 = mem_2[tmp514];
        assign tmp2024 = mem_5[tmp1950];
        assign tmp1932 = mem_2[tmp1900];
    assign tmp1898 = {temp_29[72], temp_29[73], temp_29[74], temp_29[75], temp_29[76], temp_29[77], temp_29[78], temp_29[79]};
    assign tmp2249 = tmp2247 ^ tmp2248;
    assign shifted_w3 = tmp16;
        assign tmp1556 = mem_5[tmp1489];
    assign tmp1139 = tmp1137 ^ tmp1138;
    assign tmp744 = {temp_9[104], temp_9[105], temp_9[106], temp_9[107], temp_9[108], temp_9[109], temp_9[110], temp_9[111]};
        assign tmp122 = mem_1[b2_w19];
    assign tmp2265 = tmp2263 ^ tmp2264;
        assign tmp173 = mem_1[b3_w27];
    assign b2_w31 = tmp193;
        assign tmp1841 = mem_7[tmp1725];
    assign tmp1690 = tmp1706;
        assign tmp27 = mem_3[const26_1];
    assign c4_w15 = tmp99;
    assign temp_12 = tmp953;
        assign tmp780 = mem_2[tmp748];
        assign tmp1114 = mem_6[tmp1028];
        assign tmp1314 = mem_4[tmp1255];
    assign tmp1720 = {temp_27[64], temp_27[65], temp_27[66], temp_27[67], temp_27[68], temp_27[69], temp_27[70], temp_27[71]};
        assign tmp1479 = mem_2[tmp1447];
        assign tmp1515 = mem_7[tmp1483];
    assign tmp1669 = {temp_25[64], temp_25[65], temp_25[66], temp_25[67], temp_25[68], temp_25[69], temp_25[70], temp_25[71]};
    assign tmp1816 = {tmp1815[0], tmp1815[1], tmp1815[2], tmp1815[3], tmp1815[4], tmp1815[5], tmp1815[6], tmp1815[7]};
    assign tmp1623 = tmp1621 ^ tmp1622;
    assign tmp2227 = tmp2225 ^ tmp2226;
        assign tmp2277 = mem_7[tmp2182];
    assign tmp516 = {temp_5[88], temp_5[89], temp_5[90], temp_5[91], temp_5[92], temp_5[93], temp_5[94], temp_5[95]};
    assign b1_w7 = tmp42;
    assign tmp1411 = tmp1409 ^ tmp1410;
    assign tmp25 = {c1_w3, c2_w3, c3_w3, c4_w3};
        assign tmp862 = mem_4[tmp800];
    assign tmp2111 = {temp_32[72], temp_32[73], temp_32[74], temp_32[75], temp_32[76], temp_32[77], temp_32[78], temp_32[79]};
    assign new_11 = tmp264;
        assign tmp246 = mem_1[b1_w39];
        assign tmp1239 = mem_2[tmp1207];
    assign tmp13 = {tmp11[16], tmp11[17], tmp11[18], tmp11[19], tmp11[20], tmp11[21], tmp11[22], tmp11[23]};
    assign rc3_w23 = const154_0;
    assign tmp10 = {aes_key[32], aes_key[33], aes_key[34], aes_key[35], aes_key[36], aes_key[37], aes_key[38], aes_key[39], aes_key[40], aes_key[41], aes_key[42], aes_key[43], aes_key[44], aes_key[45], aes_key[46], aes_key[47], aes_key[48], aes_key[49], aes_key[50], aes_key[51], aes_key[52], aes_key[53], aes_key[54], aes_key[55], aes_key[56], aes_key[57], aes_key[58], aes_key[59], aes_key[60], aes_key[61], aes_key[62], aes_key[63]};
    assign tmp2305 = tmp2303 ^ tmp2304;
    assign tmp1692 = tmp1708;
    assign tmp750 = {temp_9[56], temp_9[57], temp_9[58], temp_9[59], temp_9[60], temp_9[61], temp_9[62], temp_9[63]};
    assign tmp1277 = tmp1356;
    assign tmp2140 = tmp2156;
    assign tmp1054 = tmp1182;
        assign tmp828 = mem_6[tmp795];
    assign tmp1803 = tmp1801 ^ tmp1802;
    assign tmp297 = {temp_1[0], temp_1[1], temp_1[2], temp_1[3], temp_1[4], temp_1[5], temp_1[6], temp_1[7]};
        assign tmp1761 = mem_7[tmp1715];
    assign tmp793 = {temp_11[120], temp_11[121], temp_11[122], temp_11[123], temp_11[124], temp_11[125], temp_11[126], temp_11[127]};
    assign tmp439 = tmp437 ^ tmp438;
    assign tmp895 = tmp893 ^ tmp894;
    assign c2_w7 = tmp47;
        assign tmp442 = mem_4[tmp341];
    assign tmp631 = tmp629 ^ tmp630;
        assign tmp1178 = mem_6[tmp1036];
    assign tmp936 = {tmp935[0], tmp935[1], tmp935[2], tmp935[3], tmp935[4], tmp935[5], tmp935[6], tmp935[7]};
    assign tmp1229 = tmp1245;
    assign tmp1913 = tmp1929;
    assign tmp1757 = tmp1755 ^ tmp1756;
    assign tmp1977 = tmp1975 ^ tmp1976;
        assign tmp1390 = mem_5[tmp1267];
    assign tmp216 = {a2_w35, a3_w35, a4_w35, a1_w35};
    assign tmp1200 = {temp_16[0], temp_16[1], temp_16[2], temp_16[3], temp_16[4], temp_16[5], temp_16[6], temp_16[7]};
    assign c4_w19 = tmp124;
    assign tmp2129 = {temp_33[64], temp_33[65], temp_33[66], temp_33[67], temp_33[68], temp_33[69], temp_33[70], temp_33[71]};
    assign rc1_w15 = tmp102;
        assign tmp317 = mem_2[tmp285];
    assign tmp1303 = tmp1301 ^ tmp1302;
    assign tmp1732 = tmp1776;
        assign tmp2158 = mem_2[tmp2126];
    assign tmp743 = {temp_9[112], temp_9[113], temp_9[114], temp_9[115], temp_9[116], temp_9[117], temp_9[118], temp_9[119]};
    assign rc1_w31 = tmp202;
        assign tmp202 = mem_3[const201_8];
        assign tmp555 = mem_2[tmp523];
    assign tmp1967 = tmp2046;
    assign tmp1482 = temp_22 ^ tmp1481;
    assign tmp261 = tmp260 ^ tmp236;
    assign tmp682 = {tmp681[0], tmp681[1], tmp681[2], tmp681[3], tmp681[4], tmp681[5], tmp681[6], tmp681[7]};
    assign rc2_w27 = const178_0;
    assign tmp2351 = {tmp2335, tmp2348, tmp2345, tmp2342, tmp2339, tmp2336, tmp2349, tmp2346, tmp2343, tmp2340, tmp2337, tmp2350, tmp2347, tmp2344, tmp2341, tmp2338};
    assign rc3_w15 = const104_0;
    assign tmp2369 = tmp2385;
    assign tmp2114 = {temp_32[48], temp_32[49], temp_32[50], temp_32[51], temp_32[52], temp_32[53], temp_32[54], temp_32[55]};
    assign tmp1917 = tmp1933;
    assign tmp1264 = {temp_19[32], temp_19[33], temp_19[34], temp_19[35], temp_19[36], temp_19[37], temp_19[38], temp_19[39]};
        assign tmp1788 = mem_6[tmp1720];
    assign tmp1062 = {tmp1061[0], tmp1061[1], tmp1061[2], tmp1061[3], tmp1061[4], tmp1061[5], tmp1061[6], tmp1061[7]};
        assign tmp1794 = mem_5[tmp1720];
        assign tmp648 = mem_4[tmp568];
        assign tmp1801 = mem_7[tmp1720];
    assign tmp513 = {temp_5[112], temp_5[113], temp_5[114], temp_5[115], temp_5[116], temp_5[117], temp_5[118], temp_5[119]};
    assign c3_w35 = tmp223;
    assign tmp1894 = {temp_29[104], temp_29[105], temp_29[106], temp_29[107], temp_29[108], temp_29[109], temp_29[110], temp_29[111]};
    assign a3_w19 = tmp114;
    assign tmp901 = tmp899 ^ tmp900;
    assign rc4_w11 = const80_0;
    assign tmp1741 = tmp1848;
        assign tmp882 = mem_5[tmp797];
    assign tmp343 = {temp_3[40], temp_3[41], temp_3[42], temp_3[43], temp_3[44], temp_3[45], temp_3[46], temp_3[47]};
        assign tmp1298 = mem_4[tmp1253];
    assign tmp342 = {temp_3[48], temp_3[49], temp_3[50], temp_3[51], temp_3[52], temp_3[53], temp_3[54], temp_3[55]};
    assign temp_19 = new_6;
    assign tmp1530 = {tmp1529[0], tmp1529[1], tmp1529[2], tmp1529[3], tmp1529[4], tmp1529[5], tmp1529[6], tmp1529[7]};
        assign tmp1354 = mem_4[tmp1264];
    assign rc2_w15 = const103_0;
        assign tmp1928 = mem_2[tmp1896];
    assign tmp2346 = {temp_36[32], temp_36[33], temp_36[34], temp_36[35], temp_36[36], temp_36[37], temp_36[38], temp_36[39]};
        assign tmp398 = mem_5[tmp338];
    assign tmp2132 = {temp_33[40], temp_33[41], temp_33[42], temp_33[43], temp_33[44], temp_33[45], temp_33[46], temp_33[47]};
    assign tmp891 = tmp889 ^ tmp890;
        assign tmp938 = mem_5[tmp808];
    assign a2_w19 = tmp113;
        assign tmp2154 = mem_2[tmp2122];
    assign tmp2316 = {tmp2315[0], tmp2315[1], tmp2315[2], tmp2315[3], tmp2315[4], tmp2315[5], tmp2315[6], tmp2315[7]};
    assign tmp1646 = {temp_24[112], temp_24[113], temp_24[114], temp_24[115], temp_24[116], temp_24[117], temp_24[118], temp_24[119]};
    assign tmp1961 = tmp1998;
    assign tmp267 = {new_state[104], new_state[105], new_state[106], new_state[107], new_state[108], new_state[109], new_state[110], new_state[111]};
    assign tmp1807 = tmp1805 ^ tmp1806;
        assign tmp914 = mem_5[tmp801];
    assign b4_w19 = tmp120;
    assign tmp725 = {temp_8[120], temp_8[121], temp_8[122], temp_8[123], temp_8[124], temp_8[125], temp_8[126], temp_8[127]};
    assign tmp1208 = {temp_17[72], temp_17[73], temp_17[74], temp_17[75], temp_17[76], temp_17[77], temp_17[78], temp_17[79]};
        assign tmp897 = mem_7[tmp802];
    assign tmp1649 = {temp_24[88], temp_24[89], temp_24[90], temp_24[91], temp_24[92], temp_24[93], temp_24[94], temp_24[95]};
    assign tmp1412 = {tmp1411[0], tmp1411[1], tmp1411[2], tmp1411[3], tmp1411[4], tmp1411[5], tmp1411[6], tmp1411[7]};
    assign tmp1371 = tmp1369 ^ tmp1370;
        assign tmp1170 = mem_6[tmp1035];
        assign tmp1975 = mem_7[tmp1943];
        assign tmp374 = mem_5[tmp335];
    assign tmp399 = tmp397 ^ tmp398;
    assign tmp740 = {temp_8[0], temp_8[1], temp_8[2], temp_8[3], temp_8[4], temp_8[5], temp_8[6], temp_8[7]};
    assign shifted_w27 = tmp166;
    assign tmp142 = {shifted_w23[24], shifted_w23[25], shifted_w23[26], shifted_w23[27], shifted_w23[28], shifted_w23[29], shifted_w23[30], shifted_w23[31]};
    assign tmp2225 = tmp2223 ^ tmp2224;
    assign tmp1426 = {temp_20[32], temp_20[33], temp_20[34], temp_20[35], temp_20[36], temp_20[37], temp_20[38], temp_20[39]};
    assign tmp1713 = {temp_27[120], temp_27[121], temp_27[122], temp_27[123], temp_27[124], temp_27[125], temp_27[126], temp_27[127]};
    assign tmp2215 = tmp2213 ^ tmp2214;
        assign tmp1240 = mem_2[tmp1208];
    assign tmp1575 = tmp1573 ^ tmp1574;
        assign tmp1326 = mem_5[tmp1259];
        assign tmp712 = mem_4[tmp576];
    assign tmp2081 = tmp2079 ^ tmp2080;
        assign tmp1754 = mem_5[tmp1715];
    assign tmp524 = {temp_5[24], temp_5[25], temp_5[26], temp_5[27], temp_5[28], temp_5[29], temp_5[30], temp_5[31]};
    assign tmp1506 = tmp1578;
    assign tmp2038 = {tmp2037[0], tmp2037[1], tmp2037[2], tmp2037[3], tmp2037[4], tmp2037[5], tmp2037[6], tmp2037[7]};
    assign tmp657 = tmp655 ^ tmp656;
    assign tmp585 = tmp650;
        assign tmp1780 = mem_6[tmp1719];
    assign tmp1324 = {tmp1323[0], tmp1323[1], tmp1323[2], tmp1323[3], tmp1323[4], tmp1323[5], tmp1323[6], tmp1323[7]};
    assign rc1_w11 = tmp77;
    assign tmp808 = {temp_11[0], temp_11[1], temp_11[2], temp_11[3], temp_11[4], temp_11[5], temp_11[6], temp_11[7]};
    assign tmp582 = tmp626;
    assign tmp56 = {rc1_w7, rc2_w7, rc3_w7, rc4_w7};
    assign tmp2131 = {temp_33[48], temp_33[49], temp_33[50], temp_33[51], temp_33[52], temp_33[53], temp_33[54], temp_33[55]};
    assign tmp1497 = {temp_23[8], temp_23[9], temp_23[10], temp_23[11], temp_23[12], temp_23[13], temp_23[14], temp_23[15]};
    assign tmp758 = tmp774;
        assign tmp2047 = mem_7[tmp1952];
        assign tmp1534 = mem_6[tmp1483];
    assign tmp2045 = tmp2043 ^ tmp2044;
    assign tmp717 = tmp715 ^ tmp716;
    assign tmp2102 = {tmp2101[0], tmp2101[1], tmp2101[2], tmp2101[3], tmp2101[4], tmp2101[5], tmp2101[6], tmp2101[7]};
    assign tmp266 = {new_state[112], new_state[113], new_state[114], new_state[115], new_state[116], new_state[117], new_state[118], new_state[119]};
    assign b3_w31 = tmp194;
    assign tmp2352 = {temp_37[120], temp_37[121], temp_37[122], temp_37[123], temp_37[124], temp_37[125], temp_37[126], temp_37[127]};
    assign tmp2049 = tmp2047 ^ tmp2048;
        assign tmp414 = mem_5[tmp340];
        assign tmp2397 = mem_2[tmp2365];
        assign tmp1013 = mem_2[tmp981];
    assign tmp2401 = {expanded_key[1280], expanded_key[1281], expanded_key[1282], expanded_key[1283], expanded_key[1284], expanded_key[1285], expanded_key[1286], expanded_key[1287], expanded_key[1288], expanded_key[1289], expanded_key[1290], expanded_key[1291], expanded_key[1292], expanded_key[1293], expanded_key[1294], expanded_key[1295], expanded_key[1296], expanded_key[1297], expanded_key[1298], expanded_key[1299], expanded_key[1300], expanded_key[1301], expanded_key[1302], expanded_key[1303], expanded_key[1304], expanded_key[1305], expanded_key[1306], expanded_key[1307], expanded_key[1308], expanded_key[1309], expanded_key[1310], expanded_key[1311], expanded_key[1312], expanded_key[1313], expanded_key[1314], expanded_key[1315], expanded_key[1316], expanded_key[1317], expanded_key[1318], expanded_key[1319], expanded_key[1320], expanded_key[1321], expanded_key[1322], expanded_key[1323], expanded_key[1324], expanded_key[1325], expanded_key[1326], expanded_key[1327], expanded_key[1328], expanded_key[1329], expanded_key[1330], expanded_key[1331], expanded_key[1332], expanded_key[1333], expanded_key[1334], expanded_key[1335], expanded_key[1336], expanded_key[1337], expanded_key[1338], expanded_key[1339], expanded_key[1340], expanded_key[1341], expanded_key[1342], expanded_key[1343], expanded_key[1344], expanded_key[1345], expanded_key[1346], expanded_key[1347], expanded_key[1348], expanded_key[1349], expanded_key[1350], expanded_key[1351], expanded_key[1352], expanded_key[1353], expanded_key[1354], expanded_key[1355], expanded_key[1356], expanded_key[1357], expanded_key[1358], expanded_key[1359], expanded_key[1360], expanded_key[1361], expanded_key[1362], expanded_key[1363], expanded_key[1364], expanded_key[1365], expanded_key[1366], expanded_key[1367], expanded_key[1368], expanded_key[1369], expanded_key[1370], expanded_key[1371], expanded_key[1372], expanded_key[1373], expanded_key[1374], expanded_key[1375], expanded_key[1376], expanded_key[1377], expanded_key[1378], expanded_key[1379], expanded_key[1380], expanded_key[1381], expanded_key[1382], expanded_key[1383], expanded_key[1384], expanded_key[1385], expanded_key[1386], expanded_key[1387], expanded_key[1388], expanded_key[1389], expanded_key[1390], expanded_key[1391], expanded_key[1392], expanded_key[1393], expanded_key[1394], expanded_key[1395], expanded_key[1396], expanded_key[1397], expanded_key[1398], expanded_key[1399], expanded_key[1400], expanded_key[1401], expanded_key[1402], expanded_key[1403], expanded_key[1404], expanded_key[1405], expanded_key[1406], expanded_key[1407]};
    assign xor_w11 = tmp82;
    assign tmp917 = tmp915 ^ tmp916;
        assign tmp654 = mem_6[tmp568];
        assign tmp1317 = mem_7[tmp1257];
    assign temp_34 = tmp2170;
    assign shifted_w39 = tmp241;
        assign tmp1241 = mem_2[tmp1209];
    assign tmp2103 = tmp2104;
    assign tmp1227 = tmp1243;
        assign tmp1063 = mem_7[tmp1024];
        assign tmp2007 = mem_7[tmp1947];
    assign tmp1413 = tmp1414;
    assign tmp1355 = tmp1353 ^ tmp1354;
    assign tmp175 = {c1_w27, c2_w27, c3_w27, c4_w27};
    assign tmp17 = {shifted_w3[24], shifted_w3[25], shifted_w3[26], shifted_w3[27], shifted_w3[28], shifted_w3[29], shifted_w3[30], shifted_w3[31]};
        assign tmp632 = mem_4[tmp570];
    assign tmp1823 = tmp1821 ^ tmp1822;
        assign tmp2023 = mem_7[tmp1949];
    assign tmp1450 = tmp1466;
    assign tmp995 = tmp1011;
    assign tmp1840 = {tmp1839[0], tmp1839[1], tmp1839[2], tmp1839[3], tmp1839[4], tmp1839[5], tmp1839[6], tmp1839[7]};
    assign rc4_w35 = const230_0;
    assign tmp1573 = tmp1571 ^ tmp1572;
    assign tmp1907 = {temp_29[0], temp_29[1], temp_29[2], temp_29[3], temp_29[4], temp_29[5], temp_29[6], temp_29[7]};
    assign tmp1815 = tmp1813 ^ tmp1814;
    assign tmp91 = {a2_w15, a3_w15, a4_w15, a1_w15};
    assign tmp2113 = {temp_32[56], temp_32[57], temp_32[58], temp_32[59], temp_32[60], temp_32[61], temp_32[62], temp_32[63]};
    assign tmp1997 = tmp1995 ^ tmp1996;
    assign input_wire_9 = temp_6;
    assign tmp12 = {tmp11[24], tmp11[25], tmp11[26], tmp11[27], tmp11[28], tmp11[29], tmp11[30], tmp11[31]};
    assign tmp1570 = {tmp1569[0], tmp1569[1], tmp1569[2], tmp1569[3], tmp1569[4], tmp1569[5], tmp1569[6], tmp1569[7]};
    assign tmp209 = tmp208 ^ tmp184;
    assign tmp803 = {temp_11[40], temp_11[41], temp_11[42], temp_11[43], temp_11[44], temp_11[45], temp_11[46], temp_11[47]};
    assign tmp864 = {tmp863[0], tmp863[1], tmp863[2], tmp863[3], tmp863[4], tmp863[5], tmp863[6], tmp863[7]};
        assign tmp480 = mem_6[tmp345];
        assign tmp2258 = mem_4[tmp2178];
    assign tmp1843 = tmp1841 ^ tmp1842;
    assign tmp1644 = {tmp1499, tmp1500, tmp1501, tmp1502, tmp1503, tmp1504, tmp1505, tmp1506, tmp1507, tmp1508, tmp1509, tmp1510, tmp1511, tmp1512, tmp1513, tmp1514};
    assign b2_w11 = tmp68;
    assign tmp1629 = tmp1627 ^ tmp1628;
        assign tmp2240 = mem_6[tmp2179];
    assign tmp409 = tmp407 ^ tmp408;
    assign tmp361 = tmp468;
    assign tmp1545 = tmp1543 ^ tmp1544;
    assign tmp985 = {temp_13[16], temp_13[17], temp_13[18], temp_13[19], temp_13[20], temp_13[21], temp_13[22], temp_13[23]};
    assign tmp1813 = tmp1811 ^ tmp1812;
    assign tmp1853 = tmp1851 ^ tmp1852;
        assign tmp644 = mem_5[tmp570];
    assign tmp473 = tmp471 ^ tmp472;
    assign tmp745 = {temp_9[96], temp_9[97], temp_9[98], temp_9[99], temp_9[100], temp_9[101], temp_9[102], temp_9[103]};
    assign tmp411 = tmp409 ^ tmp410;
    assign tmp663 = tmp661 ^ tmp662;
        assign tmp1330 = mem_4[tmp1257];
        assign tmp1144 = mem_5[tmp1031];
        assign tmp2012 = mem_4[tmp1950];
        assign tmp552 = mem_2[tmp520];
        assign tmp249 = mem_1[b4_w39];
    assign tmp161 = tmp160 ^ tmp136;
    assign tmp1645 = {temp_24[120], temp_24[121], temp_24[122], temp_24[123], temp_24[124], temp_24[125], temp_24[126], temp_24[127]};
    assign input_wire_4 = temp_26;
    assign tmp2070 = {tmp2069[0], tmp2069[1], tmp2069[2], tmp2069[3], tmp2069[4], tmp2069[5], tmp2069[6], tmp2069[7]};
    assign tmp2356 = {temp_37[88], temp_37[89], temp_37[90], temp_37[91], temp_37[92], temp_37[93], temp_37[94], temp_37[95]};
    assign tmp731 = {temp_8[72], temp_8[73], temp_8[74], temp_8[75], temp_8[76], temp_8[77], temp_8[78], temp_8[79]};
    assign tmp1685 = tmp1701;
        assign tmp1071 = mem_7[tmp1025];
        assign tmp2387 = mem_2[tmp2355];
    assign temp_5 = tmp511;
    assign tmp331 = {expanded_key[128], expanded_key[129], expanded_key[130], expanded_key[131], expanded_key[132], expanded_key[133], expanded_key[134], expanded_key[135], expanded_key[136], expanded_key[137], expanded_key[138], expanded_key[139], expanded_key[140], expanded_key[141], expanded_key[142], expanded_key[143], expanded_key[144], expanded_key[145], expanded_key[146], expanded_key[147], expanded_key[148], expanded_key[149], expanded_key[150], expanded_key[151], expanded_key[152], expanded_key[153], expanded_key[154], expanded_key[155], expanded_key[156], expanded_key[157], expanded_key[158], expanded_key[159], expanded_key[160], expanded_key[161], expanded_key[162], expanded_key[163], expanded_key[164], expanded_key[165], expanded_key[166], expanded_key[167], expanded_key[168], expanded_key[169], expanded_key[170], expanded_key[171], expanded_key[172], expanded_key[173], expanded_key[174], expanded_key[175], expanded_key[176], expanded_key[177], expanded_key[178], expanded_key[179], expanded_key[180], expanded_key[181], expanded_key[182], expanded_key[183], expanded_key[184], expanded_key[185], expanded_key[186], expanded_key[187], expanded_key[188], expanded_key[189], expanded_key[190], expanded_key[191], expanded_key[192], expanded_key[193], expanded_key[194], expanded_key[195], expanded_key[196], expanded_key[197], expanded_key[198], expanded_key[199], expanded_key[200], expanded_key[201], expanded_key[202], expanded_key[203], expanded_key[204], expanded_key[205], expanded_key[206], expanded_key[207], expanded_key[208], expanded_key[209], expanded_key[210], expanded_key[211], expanded_key[212], expanded_key[213], expanded_key[214], expanded_key[215], expanded_key[216], expanded_key[217], expanded_key[218], expanded_key[219], expanded_key[220], expanded_key[221], expanded_key[222], expanded_key[223], expanded_key[224], expanded_key[225], expanded_key[226], expanded_key[227], expanded_key[228], expanded_key[229], expanded_key[230], expanded_key[231], expanded_key[232], expanded_key[233], expanded_key[234], expanded_key[235], expanded_key[236], expanded_key[237], expanded_key[238], expanded_key[239], expanded_key[240], expanded_key[241], expanded_key[242], expanded_key[243], expanded_key[244], expanded_key[245], expanded_key[246], expanded_key[247], expanded_key[248], expanded_key[249], expanded_key[250], expanded_key[251], expanded_key[252], expanded_key[253], expanded_key[254], expanded_key[255]};
    assign temp_32 = tmp2103;
    assign tmp754 = {temp_9[24], temp_9[25], temp_9[26], temp_9[27], temp_9[28], temp_9[29], temp_9[30], temp_9[31]};
    assign rc3_w3 = const29_0;
        assign tmp1857 = mem_7[tmp1727];
        assign tmp1017 = mem_2[tmp985];
        assign tmp1410 = mem_4[tmp1267];
        assign tmp1130 = mem_6[tmp1034];
    assign tmp330 = {tmp298, tmp299, tmp300, tmp301, tmp302, tmp303, tmp304, tmp305, tmp306, tmp307, tmp308, tmp309, tmp310, tmp311, tmp312, tmp313};
        assign tmp1098 = mem_6[tmp1030];
    assign tmp1953 = {temp_31[40], temp_31[41], temp_31[42], temp_31[43], temp_31[44], temp_31[45], temp_31[46], temp_31[47]};
        assign tmp321 = mem_2[tmp289];
    assign tmp195 = {shifted_w31[0], shifted_w31[1], shifted_w31[2], shifted_w31[3], shifted_w31[4], shifted_w31[5], shifted_w31[6], shifted_w31[7]};
        assign tmp1478 = mem_2[tmp1446];
        assign tmp2096 = mem_5[tmp1955];
    assign temp_29 = tmp1891;
        assign tmp1293 = mem_7[tmp1254];
        assign tmp1696 = mem_2[tmp1664];
        assign tmp1405 = mem_7[tmp1268];
    assign new_3 = tmp1942;
        assign tmp146 = mem_1[b1_w23];
    assign tmp2200 = tmp2300;
    assign tmp1456 = tmp1472;
    assign tmp9 = {aes_key[64], aes_key[65], aes_key[66], aes_key[67], aes_key[68], aes_key[69], aes_key[70], aes_key[71], aes_key[72], aes_key[73], aes_key[74], aes_key[75], aes_key[76], aes_key[77], aes_key[78], aes_key[79], aes_key[80], aes_key[81], aes_key[82], aes_key[83], aes_key[84], aes_key[85], aes_key[86], aes_key[87], aes_key[88], aes_key[89], aes_key[90], aes_key[91], aes_key[92], aes_key[93], aes_key[94], aes_key[95]};
    assign shifted_w31 = tmp191;
        assign tmp1978 = mem_6[tmp1945];
        assign tmp1132 = mem_4[tmp1031];
    assign tmp571 = {temp_7[56], temp_7[57], temp_7[58], temp_7[59], temp_7[60], temp_7[61], temp_7[62], temp_7[63]};
    assign tmp923 = tmp921 ^ tmp922;
    assign tmp1875 = {temp_28[120], temp_28[121], temp_28[122], temp_28[123], temp_28[124], temp_28[125], temp_28[126], temp_28[127]};
        assign tmp1938 = mem_2[tmp1906];
    assign tmp1192 = {temp_16[64], temp_16[65], temp_16[66], temp_16[67], temp_16[68], temp_16[69], temp_16[70], temp_16[71]};
        assign tmp932 = mem_6[tmp808];
        assign tmp1465 = mem_2[tmp1433];
    assign tmp278 = {new_state[16], new_state[17], new_state[18], new_state[19], new_state[20], new_state[21], new_state[22], new_state[23]};
    assign tmp1621 = tmp1619 ^ tmp1620;
        assign tmp934 = mem_4[tmp805];
    assign tmp856 = {tmp855[0], tmp855[1], tmp855[2], tmp855[3], tmp855[4], tmp855[5], tmp855[6], tmp855[7]};
    assign temp_26 = tmp1710;
    assign tmp2300 = {tmp2299[0], tmp2299[1], tmp2299[2], tmp2299[3], tmp2299[4], tmp2299[5], tmp2299[6], tmp2299[7]};
    assign tmp2195 = tmp2260;
    assign tmp1712 = temp_26 ^ tmp1711;
    assign tmp70 = {shifted_w11[0], shifted_w11[1], shifted_w11[2], shifted_w11[3], shifted_w11[4], shifted_w11[5], shifted_w11[6], shifted_w11[7]};
    assign c1_w3 = tmp21;
    assign tmp2247 = tmp2245 ^ tmp2246;
    assign tmp90 = {tmp86[0], tmp86[1], tmp86[2], tmp86[3], tmp86[4], tmp86[5], tmp86[6], tmp86[7]};
    assign tmp1527 = tmp1525 ^ tmp1526;
    assign tmp629 = tmp627 ^ tmp628;
    assign tmp653 = tmp651 ^ tmp652;
    assign tmp1969 = tmp2062;
    assign tmp1046 = tmp1118;
    assign tmp1166 = {tmp1165[0], tmp1165[1], tmp1165[2], tmp1165[3], tmp1165[4], tmp1165[5], tmp1165[6], tmp1165[7]};
    assign tmp1730 = tmp1760;
    assign tmp1213 = {temp_17[32], temp_17[33], temp_17[34], temp_17[35], temp_17[36], temp_17[37], temp_17[38], temp_17[39]};
    assign tmp2217 = tmp2215 ^ tmp2216;
        assign tmp2163 = mem_2[tmp2131];
    assign tmp1972 = tmp2086;
    assign tmp264 = aes_ciphertext ^ tmp263;
        assign tmp1167 = mem_7[tmp1037];
    assign tmp767 = tmp783;
    assign tmp62 = {tmp61[24], tmp61[25], tmp61[26], tmp61[27], tmp61[28], tmp61[29], tmp61[30], tmp61[31]};
        assign tmp2052 = mem_4[tmp1951];
        assign tmp942 = mem_4[tmp806];
        assign tmp1745 = mem_7[tmp1713];
    assign temp_24 = tmp1643;
    assign tmp277 = {new_state[24], new_state[25], new_state[26], new_state[27], new_state[28], new_state[29], new_state[30], new_state[31]};
    assign tmp1968 = tmp2054;
        assign tmp2167 = mem_2[tmp2135];
    assign tmp1952 = {temp_31[48], temp_31[49], temp_31[50], temp_31[51], temp_31[52], temp_31[53], temp_31[54], temp_31[55]};
    assign tmp133 = tmp108 ^ xor_w19;
    assign rc2_w7 = const53_0;
    assign tmp1918 = tmp1934;
    assign tmp1901 = {temp_29[48], temp_29[49], temp_29[50], temp_29[51], temp_29[52], temp_29[53], temp_29[54], temp_29[55]};
        assign tmp660 = mem_5[tmp572];
    assign tmp1270 = tmp1300;
    assign tmp641 = tmp639 ^ tmp640;
    assign c3_w19 = tmp123;
        assign tmp2386 = mem_2[tmp2354];
    assign tmp1891 = {tmp1875, tmp1888, tmp1885, tmp1882, tmp1879, tmp1876, tmp1889, tmp1886, tmp1883, tmp1880, tmp1877, tmp1890, tmp1887, tmp1884, tmp1881, tmp1878};
    assign tmp802 = {temp_11[48], temp_11[49], temp_11[50], temp_11[51], temp_11[52], temp_11[53], temp_11[54], temp_11[55]};
    assign tmp2357 = {temp_37[80], temp_37[81], temp_37[82], temp_37[83], temp_37[84], temp_37[85], temp_37[86], temp_37[87]};
    assign tmp2003 = tmp2001 ^ tmp2002;
    assign tmp508 = {temp_4[16], temp_4[17], temp_4[18], temp_4[19], temp_4[20], temp_4[21], temp_4[22], temp_4[23]};
    assign tmp2204 = tmp2332;
        assign tmp2063 = mem_7[tmp1954];
        assign tmp1074 = mem_6[tmp1023];
    assign tmp1437 = {temp_21[80], temp_21[81], temp_21[82], temp_21[83], temp_21[84], temp_21[85], temp_21[86], temp_21[87]};
    assign tmp493 = tmp494;
    assign tmp2366 = {temp_37[8], temp_37[9], temp_37[10], temp_37[11], temp_37[12], temp_37[13], temp_37[14], temp_37[15]};
        assign tmp1927 = mem_2[tmp1895];
    assign a4_w15 = tmp90;
    assign tmp1871 = tmp1869 ^ tmp1870;
    assign tmp93 = {shifted_w15[16], shifted_w15[17], shifted_w15[18], shifted_w15[19], shifted_w15[20], shifted_w15[21], shifted_w15[22], shifted_w15[23]};
    assign tmp765 = tmp781;
    assign temp_21 = tmp1431;
        assign tmp1103 = mem_7[tmp1029];
    assign a2_w15 = tmp88;
    assign tmp465 = tmp463 ^ tmp464;
        assign tmp1334 = mem_5[tmp1260];
    assign tmp510 = {temp_4[0], temp_4[1], temp_4[2], temp_4[3], temp_4[4], temp_4[5], temp_4[6], temp_4[7]};
    assign input_wire_11 = aes_ciphertext;
    assign tmp1449 = tmp1465;
        assign tmp1802 = mem_5[tmp1717];
        assign tmp370 = mem_4[tmp336];
        assign tmp1540 = mem_5[tmp1483];
        assign tmp1350 = mem_5[tmp1262];
        assign tmp1108 = mem_4[tmp1028];
        assign tmp1708 = mem_2[tmp1676];
    assign tmp1514 = tmp1642;
        assign tmp177 = mem_3[const176_7];
    assign tmp1125 = tmp1123 ^ tmp1124;
    assign tmp1666 = {temp_25[88], temp_25[89], temp_25[90], temp_25[91], temp_25[92], temp_25[93], temp_25[94], temp_25[95]};
    assign tmp1269 = tmp1292;
    assign tmp1253 = {temp_19[120], temp_19[121], temp_19[122], temp_19[123], temp_19[124], temp_19[125], temp_19[126], temp_19[127]};
    assign tmp94 = {shifted_w15[8], shifted_w15[9], shifted_w15[10], shifted_w15[11], shifted_w15[12], shifted_w15[13], shifted_w15[14], shifted_w15[15]};
    assign tmp35 = tmp34 ^ tmp10;
    assign tmp286 = {temp_1[88], temp_1[89], temp_1[90], temp_1[91], temp_1[92], temp_1[93], temp_1[94], temp_1[95]};
    assign tmp18 = {shifted_w3[16], shifted_w3[17], shifted_w3[18], shifted_w3[19], shifted_w3[20], shifted_w3[21], shifted_w3[22], shifted_w3[23]};
    assign temp_33 = tmp2121;
        assign tmp913 = mem_7[tmp804];
        assign tmp1924 = mem_2[tmp1892];
    assign tmp503 = {temp_4[56], temp_4[57], temp_4[58], temp_4[59], temp_4[60], temp_4[61], temp_4[62], temp_4[63]};
        assign tmp373 = mem_7[tmp334];
        assign tmp1774 = mem_4[tmp1715];
        assign tmp606 = mem_6[tmp566];
    assign tmp590 = tmp690;
        assign tmp638 = mem_6[tmp570];
    assign tmp335 = {temp_3[104], temp_3[105], temp_3[106], temp_3[107], temp_3[108], temp_3[109], temp_3[110], temp_3[111]};
    assign tmp1036 = {temp_15[16], temp_15[17], temp_15[18], temp_15[19], temp_15[20], temp_15[21], temp_15[22], temp_15[23]};
    assign tmp2005 = tmp2003 ^ tmp2004;
    assign tmp239 = {tmp236[8], tmp236[9], tmp236[10], tmp236[11], tmp236[12], tmp236[13], tmp236[14], tmp236[15]};
        assign tmp1234 = mem_2[tmp1202];
        assign tmp1136 = mem_5[tmp1034];
        assign tmp47 = mem_1[b2_w7];
        assign tmp2028 = mem_4[tmp1948];
    assign tmp193 = {shifted_w31[16], shifted_w31[17], shifted_w31[18], shifted_w31[19], shifted_w31[20], shifted_w31[21], shifted_w31[22], shifted_w31[23]};
    assign tmp2085 = tmp2083 ^ tmp2084;
    assign tmp1998 = {tmp1997[0], tmp1997[1], tmp1997[2], tmp1997[3], tmp1997[4], tmp1997[5], tmp1997[6], tmp1997[7]};
    assign tmp1282 = tmp1396;
    assign tmp791 = {expanded_key[384], expanded_key[385], expanded_key[386], expanded_key[387], expanded_key[388], expanded_key[389], expanded_key[390], expanded_key[391], expanded_key[392], expanded_key[393], expanded_key[394], expanded_key[395], expanded_key[396], expanded_key[397], expanded_key[398], expanded_key[399], expanded_key[400], expanded_key[401], expanded_key[402], expanded_key[403], expanded_key[404], expanded_key[405], expanded_key[406], expanded_key[407], expanded_key[408], expanded_key[409], expanded_key[410], expanded_key[411], expanded_key[412], expanded_key[413], expanded_key[414], expanded_key[415], expanded_key[416], expanded_key[417], expanded_key[418], expanded_key[419], expanded_key[420], expanded_key[421], expanded_key[422], expanded_key[423], expanded_key[424], expanded_key[425], expanded_key[426], expanded_key[427], expanded_key[428], expanded_key[429], expanded_key[430], expanded_key[431], expanded_key[432], expanded_key[433], expanded_key[434], expanded_key[435], expanded_key[436], expanded_key[437], expanded_key[438], expanded_key[439], expanded_key[440], expanded_key[441], expanded_key[442], expanded_key[443], expanded_key[444], expanded_key[445], expanded_key[446], expanded_key[447], expanded_key[448], expanded_key[449], expanded_key[450], expanded_key[451], expanded_key[452], expanded_key[453], expanded_key[454], expanded_key[455], expanded_key[456], expanded_key[457], expanded_key[458], expanded_key[459], expanded_key[460], expanded_key[461], expanded_key[462], expanded_key[463], expanded_key[464], expanded_key[465], expanded_key[466], expanded_key[467], expanded_key[468], expanded_key[469], expanded_key[470], expanded_key[471], expanded_key[472], expanded_key[473], expanded_key[474], expanded_key[475], expanded_key[476], expanded_key[477], expanded_key[478], expanded_key[479], expanded_key[480], expanded_key[481], expanded_key[482], expanded_key[483], expanded_key[484], expanded_key[485], expanded_key[486], expanded_key[487], expanded_key[488], expanded_key[489], expanded_key[490], expanded_key[491], expanded_key[492], expanded_key[493], expanded_key[494], expanded_key[495], expanded_key[496], expanded_key[497], expanded_key[498], expanded_key[499], expanded_key[500], expanded_key[501], expanded_key[502], expanded_key[503], expanded_key[504], expanded_key[505], expanded_key[506], expanded_key[507], expanded_key[508], expanded_key[509], expanded_key[510], expanded_key[511]};
        assign tmp458 = mem_4[tmp343];
    assign tmp958 = {temp_12[96], temp_12[97], temp_12[98], temp_12[99], temp_12[100], temp_12[101], temp_12[102], temp_12[103]};
        assign tmp1301 = mem_7[tmp1255];
        assign tmp1778 = mem_5[tmp1718];
    assign tmp1656 = {temp_24[32], temp_24[33], temp_24[34], temp_24[35], temp_24[36], temp_24[37], temp_24[38], temp_24[39]};
    assign tmp452 = {tmp451[0], tmp451[1], tmp451[2], tmp451[3], tmp451[4], tmp451[5], tmp451[6], tmp451[7]};
        assign tmp445 = mem_7[tmp343];
    assign tmp1903 = {temp_29[32], temp_29[33], temp_29[34], temp_29[35], temp_29[36], temp_29[37], temp_29[38], temp_29[39]};
    assign tmp1663 = {temp_25[112], temp_25[113], temp_25[114], temp_25[115], temp_25[116], temp_25[117], temp_25[118], temp_25[119]};
    assign tmp1618 = {tmp1617[0], tmp1617[1], tmp1617[2], tmp1617[3], tmp1617[4], tmp1617[5], tmp1617[6], tmp1617[7]};
    assign tmp2235 = tmp2233 ^ tmp2234;
    assign tmp1027 = {temp_15[88], temp_15[89], temp_15[90], temp_15[91], temp_15[92], temp_15[93], temp_15[94], temp_15[95]};
    assign tmp1963 = tmp2014;
    assign a1_w23 = tmp137;
    assign tmp2035 = tmp2033 ^ tmp2034;
    assign c2_w15 = tmp97;
    assign tmp2001 = tmp1999 ^ tmp2000;
    assign tmp31 = {rc1_w3, rc2_w3, rc3_w3, rc4_w3};
    assign tmp150 = {c1_w23, c2_w23, c3_w23, c4_w23};
    assign tmp282 = {temp_1[120], temp_1[121], temp_1[122], temp_1[123], temp_1[124], temp_1[125], temp_1[126], temp_1[127]};
    assign tmp407 = tmp405 ^ tmp406;
    assign tmp1053 = tmp1174;
    assign tmp1191 = {temp_16[72], temp_16[73], temp_16[74], temp_16[75], temp_16[76], temp_16[77], temp_16[78], temp_16[79]};
    assign c1_w27 = tmp171;
    assign tmp1581 = tmp1579 ^ tmp1580;
    assign input_wire_1 = temp_38;
    assign tmp132 = concat_w19 ^ substituted_w19;
    assign tmp140 = {tmp136[0], tmp136[1], tmp136[2], tmp136[3], tmp136[4], tmp136[5], tmp136[6], tmp136[7]};
    assign tmp1419 = {temp_20[88], temp_20[89], temp_20[90], temp_20[91], temp_20[92], temp_20[93], temp_20[94], temp_20[95]};
    assign tmp1323 = tmp1321 ^ tmp1322;
        assign tmp2002 = mem_6[tmp1944];
    assign shifted_w23 = tmp141;
    assign tmp1289 = tmp1287 ^ tmp1288;
    assign tmp560 = {tmp528, tmp529, tmp530, tmp531, tmp532, tmp533, tmp534, tmp535, tmp536, tmp537, tmp538, tmp539, tmp540, tmp541, tmp542, tmp543};
        assign tmp472 = mem_6[tmp348];
    assign tmp1340 = {tmp1339[0], tmp1339[1], tmp1339[2], tmp1339[3], tmp1339[4], tmp1339[5], tmp1339[6], tmp1339[7]};
    assign tmp1609 = tmp1607 ^ tmp1608;
        assign tmp2090 = mem_6[tmp1955];
        assign tmp1322 = mem_4[tmp1260];
        assign tmp884 = mem_6[tmp798];
    assign tmp1725 = {temp_27[24], temp_27[25], temp_27[26], temp_27[27], temp_27[28], temp_27[29], temp_27[30], temp_27[31]};
    assign substituted_w7 = tmp50;
    assign tmp2073 = tmp2071 ^ tmp2072;
        assign tmp1090 = mem_6[tmp1029];
        assign tmp450 = mem_4[tmp342];
    assign tmp412 = {tmp411[0], tmp411[1], tmp411[2], tmp411[3], tmp411[4], tmp411[5], tmp411[6], tmp411[7]};
    assign tmp1089 = tmp1087 ^ tmp1088;
    assign tmp1321 = tmp1319 ^ tmp1320;
        assign tmp1937 = mem_2[tmp1905];
        assign tmp2226 = mem_4[tmp2174];
        assign tmp1929 = mem_2[tmp1897];
    assign tmp1020 = {tmp988, tmp989, tmp990, tmp991, tmp992, tmp993, tmp994, tmp995, tmp996, tmp997, tmp998, tmp999, tmp1000, tmp1001, tmp1002, tmp1003};
        assign tmp397 = mem_7[tmp337];
        assign tmp1007 = mem_2[tmp975];
    assign tmp192 = {shifted_w31[24], shifted_w31[25], shifted_w31[26], shifted_w31[27], shifted_w31[28], shifted_w31[29], shifted_w31[30], shifted_w31[31]};
    assign rc3_w31 = const204_0;
        assign tmp889 = mem_7[tmp801];
    assign tmp730 = {temp_8[80], temp_8[81], temp_8[82], temp_8[83], temp_8[84], temp_8[85], temp_8[86], temp_8[87]};
    assign a1_w39 = tmp237;
    assign tmp928 = {tmp927[0], tmp927[1], tmp927[2], tmp927[3], tmp927[4], tmp927[5], tmp927[6], tmp927[7]};
        assign tmp2304 = mem_6[tmp2187];
    assign tmp867 = tmp865 ^ tmp866;
        assign tmp1703 = mem_2[tmp1671];
    assign tmp822 = tmp936;
        assign tmp248 = mem_1[b3_w39];
    assign tmp341 = {temp_3[56], temp_3[57], temp_3[58], temp_3[59], temp_3[60], temp_3[61], temp_3[62], temp_3[63]};
    assign b1_w39 = tmp242;
    assign tmp1893 = {temp_29[112], temp_29[113], temp_29[114], temp_29[115], temp_29[116], temp_29[117], temp_29[118], temp_29[119]};
    assign tmp2220 = {tmp2219[0], tmp2219[1], tmp2219[2], tmp2219[3], tmp2219[4], tmp2219[5], tmp2219[6], tmp2219[7]};
    assign tmp943 = tmp941 ^ tmp942;
    assign tmp1295 = tmp1293 ^ tmp1294;
        assign tmp1628 = mem_5[tmp1498];
    assign substituted_w27 = tmp175;
    assign tmp690 = {tmp689[0], tmp689[1], tmp689[2], tmp689[3], tmp689[4], tmp689[5], tmp689[6], tmp689[7]};
    assign tmp1776 = {tmp1775[0], tmp1775[1], tmp1775[2], tmp1775[3], tmp1775[4], tmp1775[5], tmp1775[6], tmp1775[7]};
        assign tmp1087 = mem_7[tmp1027];
    assign tmp2347 = {temp_36[24], temp_36[25], temp_36[26], temp_36[27], temp_36[28], temp_36[29], temp_36[30], temp_36[31]};
        assign tmp825 = mem_7[tmp793];
    assign tmp1950 = {temp_31[64], temp_31[65], temp_31[66], temp_31[67], temp_31[68], temp_31[69], temp_31[70], temp_31[71]};
    assign tmp1165 = tmp1163 ^ tmp1164;
    assign tmp880 = {tmp879[0], tmp879[1], tmp879[2], tmp879[3], tmp879[4], tmp879[5], tmp879[6], tmp879[7]};
        assign tmp783 = mem_2[tmp751];
    assign input_wire_2 = temp_34;
    assign tmp1944 = {temp_31[112], temp_31[113], temp_31[114], temp_31[115], temp_31[116], temp_31[117], temp_31[118], temp_31[119]};
    assign tmp1738 = tmp1824;
        assign tmp400 = mem_6[tmp339];
    assign tmp144 = {shifted_w23[8], shifted_w23[9], shifted_w23[10], shifted_w23[11], shifted_w23[12], shifted_w23[13], shifted_w23[14], shifted_w23[15]};
    assign tmp1557 = tmp1555 ^ tmp1556;
    assign tmp423 = tmp421 ^ tmp422;
    assign tmp443 = tmp441 ^ tmp442;
    assign tmp291 = {temp_1[48], temp_1[49], temp_1[50], temp_1[51], temp_1[52], temp_1[53], temp_1[54], temp_1[55]};
    assign tmp1216 = {temp_17[8], temp_17[9], temp_17[10], temp_17[11], temp_17[12], temp_17[13], temp_17[14], temp_17[15]};
    assign tmp1034 = {temp_15[32], temp_15[33], temp_15[34], temp_15[35], temp_15[36], temp_15[37], temp_15[38], temp_15[39]};
        assign tmp327 = mem_2[tmp295];
    assign tmp1848 = {tmp1847[0], tmp1847[1], tmp1847[2], tmp1847[3], tmp1847[4], tmp1847[5], tmp1847[6], tmp1847[7]};
    assign tmp65 = {tmp61[0], tmp61[1], tmp61[2], tmp61[3], tmp61[4], tmp61[5], tmp61[6], tmp61[7]};
    assign tmp417 = tmp415 ^ tmp416;
    assign tmp2170 = {tmp2138, tmp2139, tmp2140, tmp2141, tmp2142, tmp2143, tmp2144, tmp2145, tmp2146, tmp2147, tmp2148, tmp2149, tmp2150, tmp2151, tmp2152, tmp2153};
    assign tmp1942 = temp_30 ^ tmp1941;
    assign tmp1201 = {tmp1185, tmp1198, tmp1195, tmp1192, tmp1189, tmp1186, tmp1199, tmp1196, tmp1193, tmp1190, tmp1187, tmp1200, tmp1197, tmp1194, tmp1191, tmp1188};
    assign tmp1847 = tmp1845 ^ tmp1846;
    assign tmp1752 = {tmp1751[0], tmp1751[1], tmp1751[2], tmp1751[3], tmp1751[4], tmp1751[5], tmp1751[6], tmp1751[7]};
    assign xor_w27 = tmp182;
    assign tmp1287 = tmp1285 ^ tmp1286;
        assign tmp1564 = mem_5[tmp1490];
    assign c3_w27 = tmp173;
        assign tmp662 = mem_6[tmp573];
    assign tmp383 = tmp381 ^ tmp382;
        assign tmp1310 = mem_5[tmp1253];
        assign tmp1576 = mem_4[tmp1489];
    assign tmp116 = {a2_w19, a3_w19, a4_w19, a1_w19};
        assign tmp368 = mem_6[tmp335];
    assign tmp792 = temp_10 ^ tmp791;
        assign tmp921 = mem_7[tmp805];
    assign tmp1372 = {tmp1371[0], tmp1371[1], tmp1371[2], tmp1371[3], tmp1371[4], tmp1371[5], tmp1371[6], tmp1371[7]};
    assign b3_w27 = tmp169;
        assign tmp2169 = mem_2[tmp2137];
        assign tmp878 = mem_4[tmp798];
    assign tmp81 = {rc1_w11, rc2_w11, rc3_w11, rc4_w11};
    assign tmp308 = tmp324;
    assign b3_w11 = tmp69;
    assign tmp1717 = {temp_27[88], temp_27[89], temp_27[90], temp_27[91], temp_27[92], temp_27[93], temp_27[94], temp_27[95]};
    assign new_6 = tmp1252;
    assign tmp674 = {tmp673[0], tmp673[1], tmp673[2], tmp673[3], tmp673[4], tmp673[5], tmp673[6], tmp673[7]};
    assign tmp697 = tmp695 ^ tmp696;
    assign tmp2116 = {temp_32[32], temp_32[33], temp_32[34], temp_32[35], temp_32[36], temp_32[37], temp_32[38], temp_32[39]};
    assign tmp1899 = {temp_29[64], temp_29[65], temp_29[66], temp_29[67], temp_29[68], temp_29[69], temp_29[70], temp_29[71]};
    assign tmp136 = tmp135 ^ tmp111;
    assign tmp907 = tmp905 ^ tmp906;
    assign tmp2123 = {temp_33[112], temp_33[113], temp_33[114], temp_33[115], temp_33[116], temp_33[117], temp_33[118], temp_33[119]};
    assign tmp1529 = tmp1527 ^ tmp1528;
    assign tmp2257 = tmp2255 ^ tmp2256;
    assign temp_23 = new_5;
        assign tmp930 = mem_5[tmp807];
    assign tmp1805 = tmp1803 ^ tmp1804;
        assign tmp2388 = mem_2[tmp2356];
    assign tmp2273 = tmp2271 ^ tmp2272;
    assign tmp935 = tmp933 ^ tmp934;
    assign tmp888 = {tmp887[0], tmp887[1], tmp887[2], tmp887[3], tmp887[4], tmp887[5], tmp887[6], tmp887[7]};
    assign tmp1327 = tmp1325 ^ tmp1326;
    assign tmp968 = {temp_12[16], temp_12[17], temp_12[18], temp_12[19], temp_12[20], temp_12[21], temp_12[22], temp_12[23]};
        assign tmp636 = mem_5[tmp569];
    assign tmp2303 = tmp2301 ^ tmp2302;
    assign temp_38 = tmp2400;
    assign tmp996 = tmp1012;
        assign tmp1769 = mem_7[tmp1716];
    assign tmp1610 = {tmp1609[0], tmp1609[1], tmp1609[2], tmp1609[3], tmp1609[4], tmp1609[5], tmp1609[6], tmp1609[7]};
    assign a1_w27 = tmp162;
        assign tmp1701 = mem_2[tmp1669];
    assign tmp1181 = tmp1179 ^ tmp1180;
        assign tmp2214 = mem_5[tmp2175];
    assign tmp250 = {c1_w39, c2_w39, c3_w39, c4_w39};
        assign tmp2238 = mem_5[tmp2178];
        assign tmp2392 = mem_2[tmp2360];
    assign tmp271 = {new_state[72], new_state[73], new_state[74], new_state[75], new_state[76], new_state[77], new_state[78], new_state[79]};
    assign tmp927 = tmp925 ^ tmp926;
    assign shifted_w35 = tmp216;
    assign temp_22 = tmp1480;
    assign tmp574 = {temp_7[32], temp_7[33], temp_7[34], temp_7[35], temp_7[36], temp_7[37], temp_7[38], temp_7[39]};
    assign temp_3 = new_10;
        assign tmp328 = mem_2[tmp296];
    assign tmp1775 = tmp1773 ^ tmp1774;
        assign tmp1580 = mem_5[tmp1492];
    assign tmp1765 = tmp1763 ^ tmp1764;
    assign tmp1919 = tmp1935;
        assign tmp486 = mem_5[tmp345];
    assign tmp233 = tmp208 ^ xor_w35;
    assign a4_w19 = tmp115;
    assign tmp1665 = {temp_25[96], temp_25[97], temp_25[98], temp_25[99], temp_25[100], temp_25[101], temp_25[102], temp_25[103]};
        assign tmp1092 = mem_4[tmp1030];
        assign tmp640 = mem_4[tmp567];
        assign tmp2159 = mem_2[tmp2127];
    assign tmp115 = {tmp111[0], tmp111[1], tmp111[2], tmp111[3], tmp111[4], tmp111[5], tmp111[6], tmp111[7]};
    assign tmp1205 = {temp_17[96], temp_17[97], temp_17[98], temp_17[99], temp_17[100], temp_17[101], temp_17[102], temp_17[103]};
    assign tmp1591 = tmp1589 ^ tmp1590;
    assign tmp2251 = tmp2249 ^ tmp2250;
        assign tmp946 = mem_5[tmp805];
    assign tmp1864 = {tmp1863[0], tmp1863[1], tmp1863[2], tmp1863[3], tmp1863[4], tmp1863[5], tmp1863[6], tmp1863[7]};
        assign tmp1402 = mem_4[tmp1266];
        assign tmp1058 = mem_6[tmp1025];
    assign c4_w11 = tmp74;
        assign tmp2264 = mem_6[tmp2178];
    assign input_wire_7 = temp_14;
    assign tmp509 = {temp_4[8], temp_4[9], temp_4[10], temp_4[11], temp_4[12], temp_4[13], temp_4[14], temp_4[15]};
    assign tmp276 = {new_state[32], new_state[33], new_state[34], new_state[35], new_state[36], new_state[37], new_state[38], new_state[39]};
    assign c1_w15 = tmp96;
        assign tmp2396 = mem_2[tmp2364];
    assign tmp1361 = tmp1359 ^ tmp1360;
        assign tmp1826 = mem_5[tmp1724];
    assign tmp2202 = tmp2316;
    assign tmp1554 = {tmp1553[0], tmp1553[1], tmp1553[2], tmp1553[3], tmp1553[4], tmp1553[5], tmp1553[6], tmp1553[7]};
        assign tmp1996 = mem_4[tmp1944];
    assign substituted_w11 = tmp75;
        assign tmp1180 = mem_4[tmp1037];
    assign tmp1490 = {temp_23[64], temp_23[65], temp_23[66], temp_23[67], temp_23[68], temp_23[69], temp_23[70], temp_23[71]};
    assign tmp899 = tmp897 ^ tmp898;
        assign tmp1010 = mem_2[tmp978];
    assign tmp2141 = tmp2157;
    assign tmp2209 = tmp2207 ^ tmp2208;
    assign tmp1710 = {tmp1678, tmp1679, tmp1680, tmp1681, tmp1682, tmp1683, tmp1684, tmp1685, tmp1686, tmp1687, tmp1688, tmp1689, tmp1690, tmp1691, tmp1692, tmp1693};
    assign tmp2139 = tmp2155;
        assign tmp1536 = mem_4[tmp1484];
    assign tmp705 = tmp703 ^ tmp704;
    assign tmp1507 = tmp1586;
    assign tmp1687 = tmp1703;
    assign tmp764 = tmp780;
        assign tmp323 = mem_2[tmp291];
    assign tmp170 = {shifted_w27[0], shifted_w27[1], shifted_w27[2], shifted_w27[3], shifted_w27[4], shifted_w27[5], shifted_w27[6], shifted_w27[7]};
        assign tmp1608 = mem_4[tmp1493];
    assign tmp564 = {temp_7[112], temp_7[113], temp_7[114], temp_7[115], temp_7[116], temp_7[117], temp_7[118], temp_7[119]};
    assign tmp2381 = tmp2397;
        assign tmp2000 = mem_5[tmp1943];
    assign b3_w35 = tmp219;
    assign a1_w35 = tmp212;
    assign tmp2379 = tmp2395;
    assign tmp736 = {temp_8[32], temp_8[33], temp_8[34], temp_8[35], temp_8[36], temp_8[37], temp_8[38], temp_8[39]};
    assign tmp1658 = {temp_24[16], temp_24[17], temp_24[18], temp_24[19], temp_24[20], temp_24[21], temp_24[22], temp_24[23]};
    assign tmp512 = {temp_5[120], temp_5[121], temp_5[122], temp_5[123], temp_5[124], temp_5[125], temp_5[126], temp_5[127]};
    assign tmp2255 = tmp2253 ^ tmp2254;
        assign tmp715 = mem_7[tmp578];
    assign tmp1714 = {temp_27[112], temp_27[113], temp_27[114], temp_27[115], temp_27[116], temp_27[117], temp_27[118], temp_27[119]};
        assign tmp2164 = mem_2[tmp2132];
    assign tmp1432 = {temp_21[120], temp_21[121], temp_21[122], temp_21[123], temp_21[124], temp_21[125], temp_21[126], temp_21[127]};
    assign tmp925 = tmp923 ^ tmp924;
        assign tmp77 = mem_3[const76_3];
    assign tmp190 = {tmp186[0], tmp186[1], tmp186[2], tmp186[3], tmp186[4], tmp186[5], tmp186[6], tmp186[7]};
    assign c2_w23 = tmp147;
    assign tmp1599 = tmp1597 ^ tmp1598;
    assign tmp1488 = {temp_23[80], temp_23[81], temp_23[82], temp_23[83], temp_23[84], temp_23[85], temp_23[86], temp_23[87]};
    assign a4_w3 = tmp15;
    assign b2_w35 = tmp218;
    assign tmp1501 = tmp1538;
        assign tmp98 = mem_1[b3_w15];
    assign tmp280 = {new_state[0], new_state[1], new_state[2], new_state[3], new_state[4], new_state[5], new_state[6], new_state[7]};
        assign tmp322 = mem_2[tmp290];
        assign tmp426 = mem_4[tmp339];
        assign tmp2246 = mem_5[tmp2179];
    assign tmp687 = tmp685 ^ tmp686;
    assign tmp1460 = tmp1476;
    assign tmp2252 = {tmp2251[0], tmp2251[1], tmp2251[2], tmp2251[3], tmp2251[4], tmp2251[5], tmp2251[6], tmp2251[7]};
    assign tmp2077 = tmp2075 ^ tmp2076;
    assign tmp2037 = tmp2035 ^ tmp2036;
    assign tmp1586 = {tmp1585[0], tmp1585[1], tmp1585[2], tmp1585[3], tmp1585[4], tmp1585[5], tmp1585[6], tmp1585[7]};
    assign tmp947 = tmp945 ^ tmp946;
        assign tmp2320 = mem_6[tmp2185];
    assign b1_w15 = tmp92;
        assign tmp316 = mem_2[tmp284];
    assign tmp2126 = {temp_33[88], temp_33[89], temp_33[90], temp_33[91], temp_33[92], temp_33[93], temp_33[94], temp_33[95]};
    assign tmp1044 = tmp1102;
    assign a4_w39 = tmp240;
    assign tmp1331 = tmp1329 ^ tmp1330;
    assign tmp2194 = tmp2252;
    assign tmp234 = tmp233 ^ tmp209;
        assign tmp1592 = mem_4[tmp1491];
    assign tmp1149 = tmp1147 ^ tmp1148;
    assign tmp459 = tmp457 ^ tmp458;
    assign tmp1260 = {temp_19[64], temp_19[65], temp_19[66], temp_19[67], temp_19[68], temp_19[69], temp_19[70], temp_19[71]};
    assign tmp1035 = {temp_15[24], temp_15[25], temp_15[26], temp_15[27], temp_15[28], temp_15[29], temp_15[30], temp_15[31]};
        assign tmp1056 = mem_5[tmp1024];
    assign b2_w3 = tmp18;
    assign tmp994 = tmp1010;
    assign tmp189 = {tmp186[8], tmp186[9], tmp186[10], tmp186[11], tmp186[12], tmp186[13], tmp186[14], tmp186[15]};
        assign tmp1520 = mem_4[tmp1486];
    assign tmp801 = {temp_11[56], temp_11[57], temp_11[58], temp_11[59], temp_11[60], temp_11[61], temp_11[62], temp_11[63]};
        assign tmp630 = mem_6[tmp569];
        assign tmp1766 = mem_4[tmp1714];
        assign tmp1084 = mem_4[tmp1025];
    assign tmp285 = {temp_1[96], temp_1[97], temp_1[98], temp_1[99], temp_1[100], temp_1[101], temp_1[102], temp_1[103]};
    assign tmp1583 = tmp1581 ^ tmp1582;
        assign tmp1620 = mem_5[tmp1497];
        assign tmp774 = mem_2[tmp742];
    assign tmp2283 = tmp2281 ^ tmp2282;
    assign tmp1613 = tmp1611 ^ tmp1612;
    assign tmp350 = tmp380;
    assign tmp183 = tmp158 ^ xor_w27;
    assign tmp939 = tmp937 ^ tmp938;
    assign tmp1155 = tmp1153 ^ tmp1154;
    assign temp_6 = tmp560;
    assign tmp1158 = {tmp1157[0], tmp1157[1], tmp1157[2], tmp1157[3], tmp1157[4], tmp1157[5], tmp1157[6], tmp1157[7]};
    assign tmp215 = {tmp211[0], tmp211[1], tmp211[2], tmp211[3], tmp211[4], tmp211[5], tmp211[6], tmp211[7]};
    assign tmp1744 = tmp1872;
    assign tmp2021 = tmp2019 ^ tmp2020;
    assign tmp292 = {temp_1[40], temp_1[41], temp_1[42], temp_1[43], temp_1[44], temp_1[45], temp_1[46], temp_1[47]};
    assign tmp69 = {shifted_w11[8], shifted_w11[9], shifted_w11[10], shifted_w11[11], shifted_w11[12], shifted_w11[13], shifted_w11[14], shifted_w11[15]};
    assign tmp871 = tmp869 ^ tmp870;
    assign tmp1343 = tmp1341 ^ tmp1342;
    assign tmp1142 = {tmp1141[0], tmp1141[1], tmp1141[2], tmp1141[3], tmp1141[4], tmp1141[5], tmp1141[6], tmp1141[7]};
    assign tmp1956 = {temp_31[16], temp_31[17], temp_31[18], temp_31[19], temp_31[20], temp_31[21], temp_31[22], temp_31[23]};
    assign tmp597 = tmp595 ^ tmp596;
        assign tmp1096 = mem_5[tmp1029];
    assign tmp194 = {shifted_w31[8], shifted_w31[9], shifted_w31[10], shifted_w31[11], shifted_w31[12], shifted_w31[13], shifted_w31[14], shifted_w31[15]};
        assign tmp453 = mem_7[tmp344];
    assign tmp577 = {temp_7[8], temp_7[9], temp_7[10], temp_7[11], temp_7[12], temp_7[13], temp_7[14], temp_7[15]};
    assign a3_w7 = tmp39;
    assign tmp746 = {temp_9[88], temp_9[89], temp_9[90], temp_9[91], temp_9[92], temp_9[93], temp_9[94], temp_9[95]};
        assign tmp680 = mem_4[tmp572];
    assign tmp347 = {temp_3[8], temp_3[9], temp_3[10], temp_3[11], temp_3[12], temp_3[13], temp_3[14], temp_3[15]};
    assign tmp941 = tmp939 ^ tmp940;
    assign tmp2183 = {temp_35[40], temp_35[41], temp_35[42], temp_35[43], temp_35[44], temp_35[45], temp_35[46], temp_35[47]};
    assign a2_w31 = tmp188;
        assign tmp2309 = mem_7[tmp2186];
    assign tmp238 = {tmp236[16], tmp236[17], tmp236[18], tmp236[19], tmp236[20], tmp236[21], tmp236[22], tmp236[23]};
    assign tmp959 = {temp_12[88], temp_12[89], temp_12[90], temp_12[91], temp_12[92], temp_12[93], temp_12[94], temp_12[95]};
        assign tmp1309 = mem_7[tmp1256];
    assign tmp1003 = tmp1019;
    assign tmp1311 = tmp1309 ^ tmp1310;
        assign tmp1930 = mem_2[tmp1898];
        assign tmp1627 = mem_7[tmp1497];
        assign tmp97 = mem_1[b2_w15];
    assign temp_18 = tmp1250;
        assign tmp329 = mem_2[tmp297];
        assign tmp197 = mem_1[b2_w31];
    assign tmp796 = {temp_11[96], temp_11[97], temp_11[98], temp_11[99], temp_11[100], temp_11[101], temp_11[102], temp_11[103]};
    assign b4_w31 = tmp195;
        assign tmp1392 = mem_6[tmp1268];
        assign tmp198 = mem_1[b3_w31];
    assign tmp1946 = {temp_31[96], temp_31[97], temp_31[98], temp_31[99], temp_31[100], temp_31[101], temp_31[102], temp_31[103]};
        assign tmp841 = mem_7[tmp795];
    assign tmp1915 = tmp1931;
    assign tmp1308 = {tmp1307[0], tmp1307[1], tmp1307[2], tmp1307[3], tmp1307[4], tmp1307[5], tmp1307[6], tmp1307[7]};
    assign tmp58 = tmp33 ^ xor_w7;
    assign c2_w39 = tmp247;
    assign tmp1307 = tmp1305 ^ tmp1306;
        assign tmp622 = mem_6[tmp564];
        assign tmp708 = mem_5[tmp578];
    assign tmp1551 = tmp1549 ^ tmp1550;
        assign tmp1243 = mem_2[tmp1211];
    assign tmp162 = {tmp161[24], tmp161[25], tmp161[26], tmp161[27], tmp161[28], tmp161[29], tmp161[30], tmp161[31]};
    assign tmp966 = {temp_12[32], temp_12[33], temp_12[34], temp_12[35], temp_12[36], temp_12[37], temp_12[38], temp_12[39]};
    assign tmp419 = tmp417 ^ tmp418;
    assign tmp1589 = tmp1587 ^ tmp1588;
    assign tmp2287 = tmp2285 ^ tmp2286;
        assign tmp1119 = mem_7[tmp1031];
    assign tmp186 = tmp185 ^ tmp161;
        assign tmp836 = mem_6[tmp796];
    assign tmp33 = tmp8 ^ xor_w3;
        assign tmp1362 = mem_4[tmp1261];
        assign tmp1365 = mem_7[tmp1263];
        assign tmp1009 = mem_2[tmp977];
        assign tmp1707 = mem_2[tmp1675];
    assign tmp160 = tmp159 ^ tmp135;
    assign tmp1265 = {temp_19[24], temp_19[25], temp_19[26], temp_19[27], temp_19[28], temp_19[29], temp_19[30], temp_19[31]};
    assign tmp1049 = tmp1142;
    assign tmp1212 = {temp_17[40], temp_17[41], temp_17[42], temp_17[43], temp_17[44], temp_17[45], temp_17[46], temp_17[47]};
    assign tmp1693 = tmp1709;
        assign tmp2050 = mem_6[tmp1954];
    assign tmp1026 = {temp_15[96], temp_15[97], temp_15[98], temp_15[99], temp_15[100], temp_15[101], temp_15[102], temp_15[103]};
    assign input_wire_10 = temp_2;
        assign tmp777 = mem_2[tmp745];
    assign tmp455 = tmp453 ^ tmp454;
        assign tmp1563 = mem_7[tmp1489];
    assign tmp1578 = {tmp1577[0], tmp1577[1], tmp1577[2], tmp1577[3], tmp1577[4], tmp1577[5], tmp1577[6], tmp1577[7]};
    assign tmp95 = {shifted_w15[0], shifted_w15[1], shifted_w15[2], shifted_w15[3], shifted_w15[4], shifted_w15[5], shifted_w15[6], shifted_w15[7]};
        assign tmp1854 = mem_4[tmp1725];
        assign tmp2221 = mem_7[tmp2175];
        assign tmp866 = mem_5[tmp799];
        assign tmp1822 = mem_4[tmp1721];
    assign tmp1332 = {tmp1331[0], tmp1331[1], tmp1331[2], tmp1331[3], tmp1331[4], tmp1331[5], tmp1331[6], tmp1331[7]};
    assign tmp1415 = {temp_20[120], temp_20[121], temp_20[122], temp_20[123], temp_20[124], temp_20[125], temp_20[126], temp_20[127]};
    assign b4_w3 = tmp20;
    assign tmp1417 = {temp_20[104], temp_20[105], temp_20[106], temp_20[107], temp_20[108], temp_20[109], temp_20[110], temp_20[111]};
    assign tmp517 = {temp_5[80], temp_5[81], temp_5[82], temp_5[83], temp_5[84], temp_5[85], temp_5[86], temp_5[87]};
    assign tmp609 = tmp607 ^ tmp608;
    assign tmp1427 = {temp_20[24], temp_20[25], temp_20[26], temp_20[27], temp_20[28], temp_20[29], temp_20[30], temp_20[31]};
    assign tmp863 = tmp861 ^ tmp862;
        assign tmp699 = mem_7[tmp576];
    assign tmp727 = {temp_8[104], temp_8[105], temp_8[106], temp_8[107], temp_8[108], temp_8[109], temp_8[110], temp_8[111]};
        assign tmp2168 = mem_2[tmp2136];
        assign tmp1318 = mem_5[tmp1258];
    assign tmp1832 = {tmp1831[0], tmp1831[1], tmp1831[2], tmp1831[3], tmp1831[4], tmp1831[5], tmp1831[6], tmp1831[7]};
    assign b1_w31 = tmp192;
    assign tmp495 = {temp_4[120], temp_4[121], temp_4[122], temp_4[123], temp_4[124], temp_4[125], temp_4[126], temp_4[127]};
    assign a4_w23 = tmp140;
    assign tmp1727 = {temp_27[8], temp_27[9], temp_27[10], temp_27[11], temp_27[12], temp_27[13], temp_27[14], temp_27[15]};
    assign b1_w35 = tmp217;
    assign tmp1729 = tmp1752;
        assign tmp1868 = mem_6[tmp1726];
    assign tmp1498 = {temp_23[0], temp_23[1], temp_23[2], temp_23[3], temp_23[4], temp_23[5], temp_23[6], temp_23[7]};
    assign rc4_w15 = const105_0;
    assign tmp522 = {temp_5[40], temp_5[41], temp_5[42], temp_5[43], temp_5[44], temp_5[45], temp_5[46], temp_5[47]};
    assign tmp293 = {temp_1[32], temp_1[33], temp_1[34], temp_1[35], temp_1[36], temp_1[37], temp_1[38], temp_1[39]};
    assign tmp1059 = tmp1057 ^ tmp1058;
    assign tmp60 = tmp59 ^ tmp35;
    assign tmp1429 = {temp_20[8], temp_20[9], temp_20[10], temp_20[11], temp_20[12], temp_20[13], temp_20[14], temp_20[15]};
    assign tmp1233 = tmp1249;
    assign tmp358 = tmp444;
    assign tmp2135 = {temp_33[16], temp_33[17], temp_33[18], temp_33[19], temp_33[20], temp_33[21], temp_33[22], temp_33[23]};
        assign tmp1011 = mem_2[tmp979];
    assign tmp1491 = {temp_23[56], temp_23[57], temp_23[58], temp_23[59], temp_23[60], temp_23[61], temp_23[62], temp_23[63]};
    assign tmp637 = tmp635 ^ tmp636;
        assign tmp2205 = mem_7[tmp2173];
    assign concat_w15 = tmp106;
    assign tmp1945 = {temp_31[104], temp_31[105], temp_31[106], temp_31[107], temp_31[108], temp_31[109], temp_31[110], temp_31[111]};
    assign tmp1313 = tmp1311 ^ tmp1312;
    assign tmp2342 = {temp_36[64], temp_36[65], temp_36[66], temp_36[67], temp_36[68], temp_36[69], temp_36[70], temp_36[71]};
    assign b3_w15 = tmp94;
    assign tmp986 = {temp_13[8], temp_13[9], temp_13[10], temp_13[11], temp_13[12], temp_13[13], temp_13[14], temp_13[15]};
    assign tmp519 = {temp_5[64], temp_5[65], temp_5[66], temp_5[67], temp_5[68], temp_5[69], temp_5[70], temp_5[71]};
        assign tmp1175 = mem_7[tmp1038];
        assign tmp1122 = mem_6[tmp1033];
    assign tmp2029 = tmp2027 ^ tmp2028;
    assign tmp2105 = {temp_32[120], temp_32[121], temp_32[122], temp_32[123], temp_32[124], temp_32[125], temp_32[126], temp_32[127]};
        assign tmp410 = mem_4[tmp337];
    assign tmp2313 = tmp2311 ^ tmp2312;
    assign tmp1784 = {tmp1783[0], tmp1783[1], tmp1783[2], tmp1783[3], tmp1783[4], tmp1783[5], tmp1783[6], tmp1783[7]};
    assign tmp385 = tmp383 ^ tmp384;
    assign substituted_w3 = tmp25;
    assign tmp1173 = tmp1171 ^ tmp1172;
        assign tmp1064 = mem_5[tmp1025];
    assign tmp1061 = tmp1059 ^ tmp1060;
    assign tmp164 = {tmp161[8], tmp161[9], tmp161[10], tmp161[11], tmp161[12], tmp161[13], tmp161[14], tmp161[15]};
    assign tmp2236 = {tmp2235[0], tmp2235[1], tmp2235[2], tmp2235[3], tmp2235[4], tmp2235[5], tmp2235[6], tmp2235[7]};
    assign tmp496 = {temp_4[112], temp_4[113], temp_4[114], temp_4[115], temp_4[116], temp_4[117], temp_4[118], temp_4[119]};
    assign tmp1990 = {tmp1989[0], tmp1989[1], tmp1989[2], tmp1989[3], tmp1989[4], tmp1989[5], tmp1989[6], tmp1989[7]};
        assign tmp1762 = mem_5[tmp1716];
        assign tmp1830 = mem_4[tmp1722];
    assign tmp38 = {tmp36[16], tmp36[17], tmp36[18], tmp36[19], tmp36[20], tmp36[21], tmp36[22], tmp36[23]};
    assign tmp1751 = tmp1749 ^ tmp1750;
        assign tmp1247 = mem_2[tmp1215];
        assign tmp1544 = mem_4[tmp1485];
    assign b2_w39 = tmp243;
        assign tmp788 = mem_2[tmp756];
    assign tmp1086 = {tmp1085[0], tmp1085[1], tmp1085[2], tmp1085[3], tmp1085[4], tmp1085[5], tmp1085[6], tmp1085[7]};
        assign tmp1820 = mem_6[tmp1724];
    assign tmp1811 = tmp1809 ^ tmp1810;
    assign tmp1522 = {tmp1521[0], tmp1521[1], tmp1521[2], tmp1521[3], tmp1521[4], tmp1521[5], tmp1521[6], tmp1521[7]};
        assign tmp124 = mem_1[b4_w19];
        assign tmp1524 = mem_5[tmp1485];
        assign tmp614 = mem_6[tmp563];
        assign tmp1104 = mem_5[tmp1030];
    assign input_wire_8 = temp_10;
        assign tmp2095 = mem_7[tmp1958];
        assign tmp2322 = mem_4[tmp2186];
        assign tmp1082 = mem_6[tmp1024];
    assign tmp19 = {shifted_w3[8], shifted_w3[9], shifted_w3[10], shifted_w3[11], shifted_w3[12], shifted_w3[13], shifted_w3[14], shifted_w3[15]};
    assign tmp1509 = tmp1602;
        assign tmp1162 = mem_6[tmp1038];
    assign tmp1081 = tmp1079 ^ tmp1080;
    assign tmp237 = {tmp236[24], tmp236[25], tmp236[26], tmp236[27], tmp236[28], tmp236[29], tmp236[30], tmp236[31]};
    assign tmp610 = {tmp609[0], tmp609[1], tmp609[2], tmp609[3], tmp609[4], tmp609[5], tmp609[6], tmp609[7]};
    assign tmp1533 = tmp1531 ^ tmp1532;
        assign tmp1312 = mem_6[tmp1254];
    assign tmp576 = {temp_7[16], temp_7[17], temp_7[18], temp_7[19], temp_7[20], temp_7[21], temp_7[22], temp_7[23]};
    assign tmp1911 = tmp1927;
    assign tmp109 = tmp108 ^ tmp84;
    assign tmp2358 = {temp_37[72], temp_37[73], temp_37[74], temp_37[75], temp_37[76], temp_37[77], temp_37[78], temp_37[79]};
    assign tmp1032 = {temp_15[48], temp_15[49], temp_15[50], temp_15[51], temp_15[52], temp_15[53], temp_15[54], temp_15[55]};
        assign tmp704 = mem_4[tmp575];
        assign tmp2230 = mem_5[tmp2173];
    assign tmp2239 = tmp2237 ^ tmp2238;
    assign temp_27 = new_4;
        assign tmp1079 = mem_7[tmp1026];
    assign tmp1722 = {temp_27[48], temp_27[49], temp_27[50], temp_27[51], temp_27[52], temp_27[53], temp_27[54], temp_27[55]};
    assign tmp1485 = {temp_23[104], temp_23[105], temp_23[106], temp_23[107], temp_23[108], temp_23[109], temp_23[110], temp_23[111]};
        assign tmp416 = mem_6[tmp337];
    assign tmp1458 = tmp1474;
    assign tmp1031 = {temp_15[56], temp_15[57], temp_15[58], temp_15[59], temp_15[60], temp_15[61], temp_15[62], temp_15[63]};
    assign rc4_w39 = const255_0;
    assign a4_w27 = tmp165;
        assign tmp1248 = mem_2[tmp1216];
    assign tmp295 = {temp_1[16], temp_1[17], temp_1[18], temp_1[19], temp_1[20], temp_1[21], temp_1[22], temp_1[23]};
    assign tmp2137 = {temp_33[0], temp_33[1], temp_33[2], temp_33[3], temp_33[4], temp_33[5], temp_33[6], temp_33[7]};
    assign tmp1657 = {temp_24[24], temp_24[25], temp_24[26], temp_24[27], temp_24[28], temp_24[29], temp_24[30], temp_24[31]};
    assign tmp1987 = tmp1985 ^ tmp1986;
    assign tmp960 = {temp_12[80], temp_12[81], temp_12[82], temp_12[83], temp_12[84], temp_12[85], temp_12[86], temp_12[87]};
        assign tmp1936 = mem_2[tmp1904];
    assign tmp1262 = {temp_19[48], temp_19[49], temp_19[50], temp_19[51], temp_19[52], temp_19[53], temp_19[54], temp_19[55]};
    assign tmp2315 = tmp2313 ^ tmp2314;
    assign tmp1512 = tmp1626;
    assign tmp1220 = tmp1236;
    assign tmp1947 = {temp_31[88], temp_31[89], temp_31[90], temp_31[91], temp_31[92], temp_31[93], temp_31[94], temp_31[95]};
    assign b2_w15 = tmp93;
        assign tmp2222 = mem_5[tmp2176];
    assign a3_w15 = tmp89;
    assign tmp728 = {temp_8[96], temp_8[97], temp_8[98], temp_8[99], temp_8[100], temp_8[101], temp_8[102], temp_8[103]};
    assign b2_w27 = tmp168;
    assign tmp869 = tmp867 ^ tmp868;
        assign tmp2079 = mem_7[tmp1956];
    assign tmp618 = {tmp617[0], tmp617[1], tmp617[2], tmp617[3], tmp617[4], tmp617[5], tmp617[6], tmp617[7]};
    assign tmp589 = tmp682;
        assign tmp1539 = mem_7[tmp1486];
    assign tmp460 = {tmp459[0], tmp459[1], tmp459[2], tmp459[3], tmp459[4], tmp459[5], tmp459[6], tmp459[7]};
    assign tmp2184 = {temp_35[32], temp_35[33], temp_35[34], temp_35[35], temp_35[36], temp_35[37], temp_35[38], temp_35[39]};
    assign tmp1435 = {temp_21[96], temp_21[97], temp_21[98], temp_21[99], temp_21[100], temp_21[101], temp_21[102], temp_21[103]};
    assign b3_w19 = tmp119;
    assign tmp1043 = tmp1094;
    assign tmp2091 = tmp2089 ^ tmp2090;
    assign tmp1118 = {tmp1117[0], tmp1117[1], tmp1117[2], tmp1117[3], tmp1117[4], tmp1117[5], tmp1117[6], tmp1117[7]};
    assign tmp364 = tmp492;
        assign tmp366 = mem_5[tmp334];
    assign tmp580 = tmp610;
        assign tmp1603 = mem_7[tmp1494];
    assign tmp2336 = {temp_36[112], temp_36[113], temp_36[114], temp_36[115], temp_36[116], temp_36[117], temp_36[118], temp_36[119]};
    assign tmp1677 = {temp_25[0], temp_25[1], temp_25[2], temp_25[3], temp_25[4], temp_25[5], temp_25[6], temp_25[7]};
    assign tmp2299 = tmp2297 ^ tmp2298;
    assign tmp521 = {temp_5[48], temp_5[49], temp_5[50], temp_5[51], temp_5[52], temp_5[53], temp_5[54], temp_5[55]};
    assign tmp2199 = tmp2292;
        assign tmp1632 = mem_4[tmp1496];
        assign tmp2270 = mem_5[tmp2182];
    assign tmp570 = {temp_7[64], temp_7[65], temp_7[66], temp_7[67], temp_7[68], temp_7[69], temp_7[70], temp_7[71]};
        assign tmp1528 = mem_4[tmp1483];
    assign tmp1299 = tmp1297 ^ tmp1298;
    assign a3_w35 = tmp214;
        assign tmp2278 = mem_5[tmp2183];
    assign tmp588 = tmp674;
    assign tmp1923 = tmp1939;
    assign tmp1867 = tmp1865 ^ tmp1866;
    assign tmp2297 = tmp2295 ^ tmp2296;
    assign tmp967 = {temp_12[24], temp_12[25], temp_12[26], temp_12[27], temp_12[28], temp_12[29], temp_12[30], temp_12[31]};
    assign tmp1184 = {tmp1039, tmp1040, tmp1041, tmp1042, tmp1043, tmp1044, tmp1045, tmp1046, tmp1047, tmp1048, tmp1049, tmp1050, tmp1051, tmp1052, tmp1053, tmp1054};
    assign tmp2373 = tmp2389;
        assign tmp221 = mem_1[b1_w35];
        assign tmp868 = mem_6[tmp800];
    assign rc4_w31 = const205_0;
    assign tmp355 = tmp420;
        assign tmp1397 = mem_7[tmp1267];
        assign tmp1992 = mem_5[tmp1946];
    assign tmp211 = tmp210 ^ tmp186;
        assign tmp1389 = mem_7[tmp1266];
    assign c4_w35 = tmp224;
    assign tmp106 = {rc1_w15, rc2_w15, rc3_w15, rc4_w15};
    assign tmp1131 = tmp1129 ^ tmp1130;
        assign tmp860 = mem_6[tmp799];
        assign tmp1088 = mem_5[tmp1028];
    assign tmp309 = tmp325;
    assign tmp904 = {tmp903[0], tmp903[1], tmp903[2], tmp903[3], tmp903[4], tmp903[5], tmp903[6], tmp903[7]};
    assign tmp733 = {temp_8[56], temp_8[57], temp_8[58], temp_8[59], temp_8[60], temp_8[61], temp_8[62], temp_8[63]};
    assign tmp2275 = tmp2273 ^ tmp2274;
    assign tmp2011 = tmp2009 ^ tmp2010;
        assign tmp1579 = mem_7[tmp1491];
    assign tmp726 = {temp_8[112], temp_8[113], temp_8[114], temp_8[115], temp_8[116], temp_8[117], temp_8[118], temp_8[119]};
        assign tmp123 = mem_1[b3_w19];
        assign tmp2165 = mem_2[tmp2133];
    assign tmp45 = {shifted_w7[0], shifted_w7[1], shifted_w7[2], shifted_w7[3], shifted_w7[4], shifted_w7[5], shifted_w7[6], shifted_w7[7]};
    assign tmp337 = {temp_3[88], temp_3[89], temp_3[90], temp_3[91], temp_3[92], temp_3[93], temp_3[94], temp_3[95]};
    assign tmp188 = {tmp186[16], tmp186[17], tmp186[18], tmp186[19], tmp186[20], tmp186[21], tmp186[22], tmp186[23]};
    assign tmp1353 = tmp1351 ^ tmp1352;
    assign substituted_w35 = tmp225;
        assign tmp1587 = mem_7[tmp1492];
    assign b4_w11 = tmp70;
    assign tmp1549 = tmp1547 ^ tmp1548;
    assign tmp2377 = tmp2393;
    assign tmp1414 = {tmp1269, tmp1270, tmp1271, tmp1272, tmp1273, tmp1274, tmp1275, tmp1276, tmp1277, tmp1278, tmp1279, tmp1280, tmp1281, tmp1282, tmp1283, tmp1284};
    assign tmp961 = {temp_12[72], temp_12[73], temp_12[74], temp_12[75], temp_12[76], temp_12[77], temp_12[78], temp_12[79]};
    assign concat_w27 = tmp181;
    assign rc2_w11 = const78_0;
        assign tmp858 = mem_5[tmp798];
    assign c3_w3 = tmp23;
        assign tmp174 = mem_1[b4_w27];
    assign tmp1845 = tmp1843 ^ tmp1844;
    assign tmp1682 = tmp1698;
    assign tmp2371 = tmp2387;
        assign tmp1705 = mem_2[tmp1673];
    assign tmp362 = tmp476;
    assign tmp360 = tmp460;
    assign tmp1452 = tmp1468;
    assign tmp1601 = tmp1599 ^ tmp1600;
        assign tmp1552 = mem_4[tmp1490];
        assign tmp1698 = mem_2[tmp1666];
    assign tmp1163 = tmp1161 ^ tmp1162;
        assign tmp1106 = mem_6[tmp1027];
        assign tmp2084 = mem_4[tmp1955];
    assign tmp2359 = {temp_37[64], temp_37[65], temp_37[66], temp_37[67], temp_37[68], temp_37[69], temp_37[70], temp_37[71]};
    assign tmp257 = concat_w39 ^ substituted_w39;
    assign tmp1281 = tmp1388;
        assign tmp694 = mem_6[tmp577];
    assign tmp649 = tmp647 ^ tmp648;
    assign tmp1422 = {temp_20[64], temp_20[65], temp_20[66], temp_20[67], temp_20[68], temp_20[69], temp_20[70], temp_20[71]};
    assign tmp977 = {temp_13[80], temp_13[81], temp_13[82], temp_13[83], temp_13[84], temp_13[85], temp_13[86], temp_13[87]};
    assign tmp1069 = tmp1067 ^ tmp1068;
    assign tmp1424 = {temp_20[48], temp_20[49], temp_20[50], temp_20[51], temp_20[52], temp_20[53], temp_20[54], temp_20[55]};
    assign tmp877 = tmp875 ^ tmp876;
    assign tmp1487 = {temp_23[88], temp_23[89], temp_23[90], temp_23[91], temp_23[92], temp_23[93], temp_23[94], temp_23[95]};
        assign tmp545 = mem_2[tmp513];
    assign tmp2014 = {tmp2013[0], tmp2013[1], tmp2013[2], tmp2013[3], tmp2013[4], tmp2013[5], tmp2013[6], tmp2013[7]};
    assign a3_w39 = tmp239;
    assign tmp2128 = {temp_33[72], temp_33[73], temp_33[74], temp_33[75], temp_33[76], temp_33[77], temp_33[78], temp_33[79]};
    assign expanded_key = tmp262;
        assign tmp874 = mem_5[tmp800];
    assign tmp2193 = tmp2244;
    assign tmp1878 = {temp_28[96], temp_28[97], temp_28[98], temp_28[99], temp_28[100], temp_28[101], temp_28[102], temp_28[103]};
    assign temp_2 = tmp330;
    assign tmp468 = {tmp467[0], tmp467[1], tmp467[2], tmp467[3], tmp467[4], tmp467[5], tmp467[6], tmp467[7]};
        assign tmp1360 = mem_6[tmp1264];
        assign tmp2389 = mem_2[tmp2357];
        assign tmp1151 = mem_7[tmp1035];
    assign tmp498 = {temp_4[96], temp_4[97], temp_4[98], temp_4[99], temp_4[100], temp_4[101], temp_4[102], temp_4[103]};
        assign tmp2020 = mem_4[tmp1947];
        assign tmp892 = mem_6[tmp803];
    assign tmp885 = tmp883 ^ tmp884;
        assign tmp1358 = mem_5[tmp1263];
    assign tmp367 = tmp365 ^ tmp366;
    assign tmp1065 = tmp1063 ^ tmp1064;
    assign tmp1347 = tmp1345 ^ tmp1346;
        assign tmp2004 = mem_4[tmp1945];
        assign tmp1376 = mem_6[tmp1262];
    assign tmp1137 = tmp1135 ^ tmp1136;
    assign tmp1505 = tmp1570;
    assign tmp1914 = tmp1930;
    assign tmp1662 = {temp_25[120], temp_25[121], temp_25[122], temp_25[123], temp_25[124], temp_25[125], temp_25[126], temp_25[127]};
    assign tmp1940 = {tmp1908, tmp1909, tmp1910, tmp1911, tmp1912, tmp1913, tmp1914, tmp1915, tmp1916, tmp1917, tmp1918, tmp1919, tmp1920, tmp1921, tmp1922, tmp1923};
        assign tmp1068 = mem_4[tmp1023];
    assign tmp795 = {temp_11[104], temp_11[105], temp_11[106], temp_11[107], temp_11[108], temp_11[109], temp_11[110], temp_11[111]};
        assign tmp785 = mem_2[tmp753];
        assign tmp148 = mem_1[b3_w23];
    assign new_10 = tmp332;
        assign tmp1770 = mem_5[tmp1713];
    assign tmp1261 = {temp_19[56], temp_19[57], temp_19[58], temp_19[59], temp_19[60], temp_19[61], temp_19[62], temp_19[63]};
        assign tmp1014 = mem_2[tmp982];
        assign tmp779 = mem_2[tmp747];
    assign tmp2046 = {tmp2045[0], tmp2045[1], tmp2045[2], tmp2045[3], tmp2045[4], tmp2045[5], tmp2045[6], tmp2045[7]};
        assign tmp1866 = mem_5[tmp1725];
    assign tmp987 = {temp_13[0], temp_13[1], temp_13[2], temp_13[3], temp_13[4], temp_13[5], temp_13[6], temp_13[7]};
    assign tmp1920 = tmp1936;
    assign tmp1315 = tmp1313 ^ tmp1314;
    assign tmp1209 = {temp_17[64], temp_17[65], temp_17[66], temp_17[67], temp_17[68], temp_17[69], temp_17[70], temp_17[71]};
    assign tmp1225 = tmp1241;
    assign tmp1718 = {temp_27[80], temp_27[81], temp_27[82], temp_27[83], temp_27[84], temp_27[85], temp_27[86], temp_27[87]};
    assign tmp1101 = tmp1099 ^ tmp1100;
    assign tmp2069 = tmp2067 ^ tmp2068;
    assign tmp944 = {tmp943[0], tmp943[1], tmp943[2], tmp943[3], tmp943[4], tmp943[5], tmp943[6], tmp943[7]};
        assign tmp1370 = mem_4[tmp1262];
    assign tmp561 = {expanded_key[256], expanded_key[257], expanded_key[258], expanded_key[259], expanded_key[260], expanded_key[261], expanded_key[262], expanded_key[263], expanded_key[264], expanded_key[265], expanded_key[266], expanded_key[267], expanded_key[268], expanded_key[269], expanded_key[270], expanded_key[271], expanded_key[272], expanded_key[273], expanded_key[274], expanded_key[275], expanded_key[276], expanded_key[277], expanded_key[278], expanded_key[279], expanded_key[280], expanded_key[281], expanded_key[282], expanded_key[283], expanded_key[284], expanded_key[285], expanded_key[286], expanded_key[287], expanded_key[288], expanded_key[289], expanded_key[290], expanded_key[291], expanded_key[292], expanded_key[293], expanded_key[294], expanded_key[295], expanded_key[296], expanded_key[297], expanded_key[298], expanded_key[299], expanded_key[300], expanded_key[301], expanded_key[302], expanded_key[303], expanded_key[304], expanded_key[305], expanded_key[306], expanded_key[307], expanded_key[308], expanded_key[309], expanded_key[310], expanded_key[311], expanded_key[312], expanded_key[313], expanded_key[314], expanded_key[315], expanded_key[316], expanded_key[317], expanded_key[318], expanded_key[319], expanded_key[320], expanded_key[321], expanded_key[322], expanded_key[323], expanded_key[324], expanded_key[325], expanded_key[326], expanded_key[327], expanded_key[328], expanded_key[329], expanded_key[330], expanded_key[331], expanded_key[332], expanded_key[333], expanded_key[334], expanded_key[335], expanded_key[336], expanded_key[337], expanded_key[338], expanded_key[339], expanded_key[340], expanded_key[341], expanded_key[342], expanded_key[343], expanded_key[344], expanded_key[345], expanded_key[346], expanded_key[347], expanded_key[348], expanded_key[349], expanded_key[350], expanded_key[351], expanded_key[352], expanded_key[353], expanded_key[354], expanded_key[355], expanded_key[356], expanded_key[357], expanded_key[358], expanded_key[359], expanded_key[360], expanded_key[361], expanded_key[362], expanded_key[363], expanded_key[364], expanded_key[365], expanded_key[366], expanded_key[367], expanded_key[368], expanded_key[369], expanded_key[370], expanded_key[371], expanded_key[372], expanded_key[373], expanded_key[374], expanded_key[375], expanded_key[376], expanded_key[377], expanded_key[378], expanded_key[379], expanded_key[380], expanded_key[381], expanded_key[382], expanded_key[383]};
    assign tmp851 = tmp849 ^ tmp850;
    assign tmp44 = {shifted_w7[8], shifted_w7[9], shifted_w7[10], shifted_w7[11], shifted_w7[12], shifted_w7[13], shifted_w7[14], shifted_w7[15]};
    assign tmp2323 = tmp2321 ^ tmp2322;
        assign tmp252 = mem_3[const251_10];
        assign tmp2042 = mem_6[tmp1953];
    assign tmp500 = {temp_4[80], temp_4[81], temp_4[82], temp_4[83], temp_4[84], temp_4[85], temp_4[86], temp_4[87]};
        assign tmp1865 = mem_7[tmp1728];
    assign tmp82 = concat_w11 ^ substituted_w11;
    assign tmp1905 = {temp_29[16], temp_29[17], temp_29[18], temp_29[19], temp_29[20], temp_29[21], temp_29[22], temp_29[23]};
    assign tmp302 = tmp318;
        assign tmp2318 = mem_5[tmp2188];
    assign tmp167 = {shifted_w27[24], shifted_w27[25], shifted_w27[26], shifted_w27[27], shifted_w27[28], shifted_w27[29], shifted_w27[30], shifted_w27[31]};
    assign tmp489 = tmp487 ^ tmp488;
        assign tmp1357 = mem_7[tmp1262];
    assign tmp2133 = {temp_33[32], temp_33[33], temp_33[34], temp_33[35], temp_33[36], temp_33[37], temp_33[38], temp_33[39]};
    assign tmp2150 = tmp2166;
        assign tmp448 = mem_6[tmp341];
    assign tmp2374 = tmp2390;
    assign tmp806 = {temp_11[16], temp_11[17], temp_11[18], temp_11[19], temp_11[20], temp_11[21], temp_11[22], temp_11[23]};
        assign tmp2262 = mem_5[tmp2177];
    assign tmp1648 = {temp_24[96], temp_24[97], temp_24[98], temp_24[99], temp_24[100], temp_24[101], temp_24[102], temp_24[103]};
    assign tmp583 = tmp634;
    assign tmp1057 = tmp1055 ^ tmp1056;
    assign rc3_w27 = const179_0;
    assign tmp593 = tmp714;
    assign tmp100 = {c1_w15, c2_w15, c3_w15, c4_w15};
    assign tmp1492 = {temp_23[48], temp_23[49], temp_23[50], temp_23[51], temp_23[52], temp_23[53], temp_23[54], temp_23[55]};
    assign tmp1948 = {temp_31[80], temp_31[81], temp_31[82], temp_31[83], temp_31[84], temp_31[85], temp_31[86], temp_31[87]};
        assign tmp2055 = mem_7[tmp1953];
    assign b1_w19 = tmp117;
        assign tmp611 = mem_7[tmp565];
        assign tmp440 = mem_6[tmp344];
    assign tmp1675 = {temp_25[16], temp_25[17], temp_25[18], temp_25[19], temp_25[20], temp_25[21], temp_25[22], temp_25[23]};
    assign input_wire_5 = temp_22;
        assign tmp1999 = mem_7[tmp1946];
        assign tmp1246 = mem_2[tmp1214];
    assign tmp1876 = {temp_28[112], temp_28[113], temp_28[114], temp_28[115], temp_28[116], temp_28[117], temp_28[118], temp_28[119]};
    assign tmp57 = concat_w7 ^ substituted_w7;
        assign tmp1111 = mem_7[tmp1030];
    assign tmp1895 = {temp_29[96], temp_29[97], temp_29[98], temp_29[99], temp_29[100], temp_29[101], temp_29[102], temp_29[103]};
    assign tmp1067 = tmp1065 ^ tmp1066;
    assign tmp992 = tmp1008;
    assign tmp1859 = tmp1857 ^ tmp1858;
    assign tmp2051 = tmp2049 ^ tmp2050;
        assign tmp1346 = mem_4[tmp1259];
        assign tmp1571 = mem_7[tmp1490];
    assign tmp2115 = {temp_32[40], temp_32[41], temp_32[42], temp_32[43], temp_32[44], temp_32[45], temp_32[46], temp_32[47]};
    assign tmp2289 = tmp2287 ^ tmp2288;
    assign concat_w3 = tmp31;
        assign tmp466 = mem_4[tmp348];
    assign tmp2118 = {temp_32[16], temp_32[17], temp_32[18], temp_32[19], temp_32[20], temp_32[21], temp_32[22], temp_32[23]};
    assign tmp42 = {shifted_w7[24], shifted_w7[25], shifted_w7[26], shifted_w7[27], shifted_w7[28], shifted_w7[29], shifted_w7[30], shifted_w7[31]};
    assign tmp1305 = tmp1303 ^ tmp1304;
        assign tmp1931 = mem_2[tmp1899];
    assign tmp401 = tmp399 ^ tmp400;
    assign tmp1869 = tmp1867 ^ tmp1868;
        assign tmp2074 = mem_6[tmp1957];
    assign rc1_w39 = tmp252;
    assign c1_w19 = tmp121;
    assign tmp357 = tmp436;
    assign tmp642 = {tmp641[0], tmp641[1], tmp641[2], tmp641[3], tmp641[4], tmp641[5], tmp641[6], tmp641[7]};
    assign tmp605 = tmp603 ^ tmp604;
    assign tmp2259 = tmp2257 ^ tmp2258;
    assign tmp1650 = {temp_24[80], temp_24[81], temp_24[82], temp_24[83], temp_24[84], temp_24[85], temp_24[86], temp_24[87]};
    assign tmp1561 = tmp1559 ^ tmp1560;
        assign tmp1523 = mem_7[tmp1484];
        assign tmp2160 = mem_2[tmp2128];
        assign tmp2016 = mem_5[tmp1949];
    assign tmp1147 = tmp1145 ^ tmp1146;
    assign tmp2354 = {temp_37[104], temp_37[105], temp_37[106], temp_37[107], temp_37[108], temp_37[109], temp_37[110], temp_37[111]};
    assign tmp1922 = tmp1938;
    assign tmp1204 = {temp_17[104], temp_17[105], temp_17[106], temp_17[107], temp_17[108], temp_17[109], temp_17[110], temp_17[111]};
        assign tmp1135 = mem_7[tmp1033];
        assign tmp2234 = mem_4[tmp2175];
        assign tmp405 = mem_7[tmp338];
        assign tmp684 = mem_5[tmp571];
        assign tmp1984 = mem_5[tmp1945];
    assign tmp2311 = tmp2309 ^ tmp2310;
        assign tmp2071 = mem_7[tmp1955];
    assign tmp507 = {temp_4[24], temp_4[25], temp_4[26], temp_4[27], temp_4[28], temp_4[29], temp_4[30], temp_4[31]};
        assign tmp1019 = mem_2[tmp987];
    assign tmp810 = tmp840;
        assign tmp786 = mem_2[tmp754];
        assign tmp462 = mem_5[tmp346];
    assign tmp2207 = tmp2205 ^ tmp2206;
    assign tmp1489 = {temp_23[72], temp_23[73], temp_23[74], temp_23[75], temp_23[76], temp_23[77], temp_23[78], temp_23[79]};
        assign tmp852 = mem_6[tmp794];
    assign tmp467 = tmp465 ^ tmp466;
    assign c2_w19 = tmp122;
    assign tmp518 = {temp_5[72], temp_5[73], temp_5[74], temp_5[75], temp_5[76], temp_5[77], temp_5[78], temp_5[79]};
    assign tmp1569 = tmp1567 ^ tmp1568;
        assign tmp553 = mem_2[tmp521];
    assign tmp1423 = {temp_20[56], temp_20[57], temp_20[58], temp_20[59], temp_20[60], temp_20[61], temp_20[62], temp_20[63]};
    assign a3_w27 = tmp164;
    assign tmp117 = {shifted_w19[24], shifted_w19[25], shifted_w19[26], shifted_w19[27], shifted_w19[28], shifted_w19[29], shifted_w19[30], shifted_w19[31]};
    assign tmp1416 = {temp_20[112], temp_20[113], temp_20[114], temp_20[115], temp_20[116], temp_20[117], temp_20[118], temp_20[119]};
    assign tmp165 = {tmp161[0], tmp161[1], tmp161[2], tmp161[3], tmp161[4], tmp161[5], tmp161[6], tmp161[7]};
        assign tmp1384 = mem_6[tmp1267];
    assign tmp953 = tmp954;
    assign tmp976 = {temp_13[88], temp_13[89], temp_13[90], temp_13[91], temp_13[92], temp_13[93], temp_13[94], temp_13[95]};
    assign tmp829 = tmp827 ^ tmp828;
        assign tmp1606 = mem_6[tmp1492];
    assign tmp112 = {tmp111[24], tmp111[25], tmp111[26], tmp111[27], tmp111[28], tmp111[29], tmp111[30], tmp111[31]};
    assign tmp1276 = tmp1348;
        assign tmp2058 = mem_6[tmp1951];
        assign tmp149 = mem_1[b4_w23];
    assign tmp584 = tmp642;
    assign tmp1486 = {temp_23[96], temp_23[97], temp_23[98], temp_23[99], temp_23[100], temp_23[101], temp_23[102], temp_23[103]};
    assign rc2_w23 = const153_0;
        assign tmp1630 = mem_6[tmp1495];
    assign tmp2043 = tmp2041 ^ tmp2042;
    assign tmp471 = tmp469 ^ tmp470;
    assign tmp1292 = {tmp1291[0], tmp1291[1], tmp1291[2], tmp1291[3], tmp1291[4], tmp1291[5], tmp1291[6], tmp1291[7]};
    assign tmp2172 = temp_34 ^ tmp2171;
    assign tmp2201 = tmp2308;
    assign tmp2223 = tmp2221 ^ tmp2222;
    assign tmp1993 = tmp1991 ^ tmp1992;
        assign tmp1986 = mem_6[tmp1946];
    assign input_wire_3 = temp_30;
        assign tmp1976 = mem_5[tmp1944];
        assign tmp850 = mem_5[tmp793];
    assign tmp428 = {tmp427[0], tmp427[1], tmp427[2], tmp427[3], tmp427[4], tmp427[5], tmp427[6], tmp427[7]};
    assign tmp1179 = tmp1177 ^ tmp1178;
    assign tmp1900 = {temp_29[56], temp_29[57], temp_29[58], temp_29[59], temp_29[60], temp_29[61], temp_29[62], temp_29[63]};
    assign tmp768 = tmp784;
    assign tmp120 = {shifted_w19[0], shifted_w19[1], shifted_w19[2], shifted_w19[3], shifted_w19[4], shifted_w19[5], shifted_w19[6], shifted_w19[7]};
    assign tmp1884 = {temp_28[48], temp_28[49], temp_28[50], temp_28[51], temp_28[52], temp_28[53], temp_28[54], temp_28[55]};
    assign tmp283 = {temp_1[112], temp_1[113], temp_1[114], temp_1[115], temp_1[116], temp_1[117], temp_1[118], temp_1[119]};
        assign tmp2301 = mem_7[tmp2185];
        assign tmp1100 = mem_4[tmp1027];
        assign tmp2015 = mem_7[tmp1948];
    assign tmp872 = {tmp871[0], tmp871[1], tmp871[2], tmp871[3], tmp871[4], tmp871[5], tmp871[6], tmp871[7]};
    assign tmp1141 = tmp1139 ^ tmp1140;
        assign tmp1406 = mem_5[tmp1265];
    assign tmp1559 = tmp1557 ^ tmp1558;
    assign tmp2338 = {temp_36[96], temp_36[97], temp_36[98], temp_36[99], temp_36[100], temp_36[101], temp_36[102], temp_36[103]};
    assign tmp1150 = {tmp1149[0], tmp1149[1], tmp1149[2], tmp1149[3], tmp1149[4], tmp1149[5], tmp1149[6], tmp1149[7]};
    assign tmp915 = tmp913 ^ tmp914;
    assign temp_15 = new_7;
    assign tmp2125 = {temp_33[96], temp_33[97], temp_33[98], temp_33[99], temp_33[100], temp_33[101], temp_33[102], temp_33[103]};
    assign tmp1724 = {temp_27[32], temp_27[33], temp_27[34], temp_27[35], temp_27[36], temp_27[37], temp_27[38], temp_27[39]};
    assign shifted_w15 = tmp91;
        assign tmp784 = mem_2[tmp752];
    assign tmp2134 = {temp_33[24], temp_33[25], temp_33[26], temp_33[27], temp_33[28], temp_33[29], temp_33[30], temp_33[31]};
    assign tmp262 = {tmp8, tmp9, tmp10, tmp11, tmp33, tmp34, tmp35, tmp36, tmp58, tmp59, tmp60, tmp61, tmp83, tmp84, tmp85, tmp86, tmp108, tmp109, tmp110, tmp111, tmp133, tmp134, tmp135, tmp136, tmp158, tmp159, tmp160, tmp161, tmp183, tmp184, tmp185, tmp186, tmp208, tmp209, tmp210, tmp211, tmp233, tmp234, tmp235, tmp236, tmp258, tmp259, tmp260, tmp261};
    assign tmp1747 = tmp1745 ^ tmp1746;
    assign tmp820 = tmp920;
    assign new_1 = tmp2402;
    assign tmp2119 = {temp_32[8], temp_32[9], temp_32[10], temp_32[11], temp_32[12], temp_32[13], temp_32[14], temp_32[15]};
    assign xor_w39 = tmp257;
        assign tmp2229 = mem_7[tmp2176];
        assign tmp1600 = mem_4[tmp1492];
    assign tmp463 = tmp461 ^ tmp462;
        assign tmp2310 = mem_5[tmp2187];
    assign tmp729 = {temp_8[88], temp_8[89], temp_8[90], temp_8[91], temp_8[92], temp_8[93], temp_8[94], temp_8[95]};
        assign tmp2216 = mem_6[tmp2176];
    assign tmp1723 = {temp_27[40], temp_27[41], temp_27[42], temp_27[43], temp_27[44], temp_27[45], temp_27[46], temp_27[47]};
    assign tmp2122 = {temp_33[120], temp_33[121], temp_33[122], temp_33[123], temp_33[124], temp_33[125], temp_33[126], temp_33[127]};
    assign tmp1882 = {temp_28[64], temp_28[65], temp_28[66], temp_28[67], temp_28[68], temp_28[69], temp_28[70], temp_28[71]};
    assign tmp1916 = tmp1932;
    assign tmp1206 = {temp_17[88], temp_17[89], temp_17[90], temp_17[91], temp_17[92], temp_17[93], temp_17[94], temp_17[95]};
        assign tmp842 = mem_5[tmp796];
    assign xor_w7 = tmp57;
    assign concat_w7 = tmp56;
    assign tmp1194 = {temp_16[48], temp_16[49], temp_16[50], temp_16[51], temp_16[52], temp_16[53], temp_16[54], temp_16[55]};
        assign tmp1146 = mem_6[tmp1032];
    assign tmp2097 = tmp2095 ^ tmp2096;
    assign tmp235 = tmp234 ^ tmp210;
    assign tmp273 = {new_state[56], new_state[57], new_state[58], new_state[59], new_state[60], new_state[61], new_state[62], new_state[63]};
    assign tmp949 = tmp947 ^ tmp948;
        assign tmp1699 = mem_2[tmp1667];
    assign tmp1283 = tmp1404;
        assign tmp778 = mem_2[tmp746];
    assign tmp1274 = tmp1332;
    assign tmp669 = tmp667 ^ tmp668;
        assign tmp659 = mem_7[tmp571];
    assign tmp1543 = tmp1541 ^ tmp1542;
    assign tmp763 = tmp779;
        assign tmp781 = mem_2[tmp749];
    assign tmp89 = {tmp86[8], tmp86[9], tmp86[10], tmp86[11], tmp86[12], tmp86[13], tmp86[14], tmp86[15]};
    assign tmp819 = tmp912;
        assign tmp2266 = mem_4[tmp2179];
        assign tmp1472 = mem_2[tmp1440];
    assign tmp1051 = tmp1158;
    assign tmp1856 = {tmp1855[0], tmp1855[1], tmp1855[2], tmp1855[3], tmp1855[4], tmp1855[5], tmp1855[6], tmp1855[7]};
    assign tmp1827 = tmp1825 ^ tmp1826;
        assign tmp1604 = mem_5[tmp1491];
        assign tmp830 = mem_4[tmp796];
    assign tmp1428 = {temp_20[16], temp_20[17], temp_20[18], temp_20[19], temp_20[20], temp_20[21], temp_20[22], temp_20[23]};
        assign tmp924 = mem_6[tmp807];
    assign rc3_w11 = const79_0;
    assign tmp1995 = tmp1993 ^ tmp1994;
    assign tmp1639 = tmp1637 ^ tmp1638;
    assign tmp1222 = tmp1238;
    assign tmp818 = tmp904;
    assign tmp1767 = tmp1765 ^ tmp1766;
    assign tmp50 = {c1_w7, c2_w7, c3_w7, c4_w7};
    assign tmp1921 = tmp1937;
        assign tmp1304 = mem_6[tmp1253];
    assign tmp753 = {temp_9[32], temp_9[33], temp_9[34], temp_9[35], temp_9[36], temp_9[37], temp_9[38], temp_9[39]};
        assign tmp1753 = mem_7[tmp1714];
    assign tmp2182 = {temp_35[48], temp_35[49], temp_35[50], temp_35[51], temp_35[52], temp_35[53], temp_35[54], temp_35[55]};
    assign tmp1396 = {tmp1395[0], tmp1395[1], tmp1395[2], tmp1395[3], tmp1395[4], tmp1395[5], tmp1395[6], tmp1395[7]};
    assign tmp1679 = tmp1695;
    assign tmp832 = {tmp831[0], tmp831[1], tmp831[2], tmp831[3], tmp831[4], tmp831[5], tmp831[6], tmp831[7]};
    assign tmp1297 = tmp1295 ^ tmp1296;
        assign tmp2395 = mem_2[tmp2363];
        assign tmp620 = mem_5[tmp563];
        assign tmp1748 = mem_6[tmp1715];
        assign tmp1386 = mem_4[tmp1268];
    assign tmp475 = tmp473 ^ tmp474;
        assign tmp2237 = mem_7[tmp2177];
    assign tmp835 = tmp833 ^ tmp834;
    assign tmp166 = {a2_w27, a3_w27, a4_w27, a1_w27};
    assign tmp2083 = tmp2081 ^ tmp2082;
    assign tmp274 = {new_state[48], new_state[49], new_state[50], new_state[51], new_state[52], new_state[53], new_state[54], new_state[55]};
    assign tmp1835 = tmp1833 ^ tmp1834;
    assign tmp1448 = tmp1464;
    assign tmp903 = tmp901 ^ tmp902;
        assign tmp678 = mem_6[tmp571];
        assign tmp1008 = mem_2[tmp976];
        assign tmp1612 = mem_5[tmp1496];
    assign tmp817 = tmp896;
    assign rc3_w7 = const54_0;
    assign tmp219 = {shifted_w35[8], shifted_w35[9], shifted_w35[10], shifted_w35[11], shifted_w35[12], shifted_w35[13], shifted_w35[14], shifted_w35[15]};
        assign tmp1796 = mem_6[tmp1717];
    assign tmp2334 = {tmp2189, tmp2190, tmp2191, tmp2192, tmp2193, tmp2194, tmp2195, tmp2196, tmp2197, tmp2198, tmp2199, tmp2200, tmp2201, tmp2202, tmp2203, tmp2204};
        assign tmp2044 = mem_4[tmp1954];
    assign tmp1210 = {temp_17[56], temp_17[57], temp_17[58], temp_17[59], temp_17[60], temp_17[61], temp_17[62], temp_17[63]};
    assign a3_w11 = tmp64;
    assign tmp310 = tmp326;
        assign tmp905 = mem_7[tmp803];
        assign tmp1004 = mem_2[tmp972];
        assign tmp464 = mem_6[tmp347];
        assign tmp656 = mem_4[tmp569];
    assign tmp1356 = {tmp1355[0], tmp1355[1], tmp1355[2], tmp1355[3], tmp1355[4], tmp1355[5], tmp1355[6], tmp1355[7]};
        assign tmp1636 = mem_5[tmp1495];
    assign c1_w35 = tmp221;
    assign tmp2372 = tmp2388;
    assign tmp1256 = {temp_19[96], temp_19[97], temp_19[98], temp_19[99], temp_19[100], temp_19[101], temp_19[102], temp_19[103]};
    assign tmp1457 = tmp1473;
    assign temp_20 = tmp1413;
    assign tmp2268 = {tmp2267[0], tmp2267[1], tmp2267[2], tmp2267[3], tmp2267[4], tmp2267[5], tmp2267[6], tmp2267[7]};
    assign temp_30 = tmp1940;
    assign tmp535 = tmp551;
    assign tmp231 = {rc1_w35, rc2_w35, rc3_w35, rc4_w35};
    assign tmp1436 = {temp_21[88], temp_21[89], temp_21[90], temp_21[91], temp_21[92], temp_21[93], temp_21[94], temp_21[95]};
    assign tmp766 = tmp782;
        assign tmp1333 = mem_7[tmp1259];
    assign c3_w11 = tmp73;
        assign tmp1709 = mem_2[tmp1677];
    assign tmp1742 = tmp1856;
        assign tmp1790 = mem_4[tmp1717];
    assign tmp2151 = tmp2167;
    assign tmp722 = {tmp721[0], tmp721[1], tmp721[2], tmp721[3], tmp721[4], tmp721[5], tmp721[6], tmp721[7]};
    assign tmp1251 = {expanded_key[640], expanded_key[641], expanded_key[642], expanded_key[643], expanded_key[644], expanded_key[645], expanded_key[646], expanded_key[647], expanded_key[648], expanded_key[649], expanded_key[650], expanded_key[651], expanded_key[652], expanded_key[653], expanded_key[654], expanded_key[655], expanded_key[656], expanded_key[657], expanded_key[658], expanded_key[659], expanded_key[660], expanded_key[661], expanded_key[662], expanded_key[663], expanded_key[664], expanded_key[665], expanded_key[666], expanded_key[667], expanded_key[668], expanded_key[669], expanded_key[670], expanded_key[671], expanded_key[672], expanded_key[673], expanded_key[674], expanded_key[675], expanded_key[676], expanded_key[677], expanded_key[678], expanded_key[679], expanded_key[680], expanded_key[681], expanded_key[682], expanded_key[683], expanded_key[684], expanded_key[685], expanded_key[686], expanded_key[687], expanded_key[688], expanded_key[689], expanded_key[690], expanded_key[691], expanded_key[692], expanded_key[693], expanded_key[694], expanded_key[695], expanded_key[696], expanded_key[697], expanded_key[698], expanded_key[699], expanded_key[700], expanded_key[701], expanded_key[702], expanded_key[703], expanded_key[704], expanded_key[705], expanded_key[706], expanded_key[707], expanded_key[708], expanded_key[709], expanded_key[710], expanded_key[711], expanded_key[712], expanded_key[713], expanded_key[714], expanded_key[715], expanded_key[716], expanded_key[717], expanded_key[718], expanded_key[719], expanded_key[720], expanded_key[721], expanded_key[722], expanded_key[723], expanded_key[724], expanded_key[725], expanded_key[726], expanded_key[727], expanded_key[728], expanded_key[729], expanded_key[730], expanded_key[731], expanded_key[732], expanded_key[733], expanded_key[734], expanded_key[735], expanded_key[736], expanded_key[737], expanded_key[738], expanded_key[739], expanded_key[740], expanded_key[741], expanded_key[742], expanded_key[743], expanded_key[744], expanded_key[745], expanded_key[746], expanded_key[747], expanded_key[748], expanded_key[749], expanded_key[750], expanded_key[751], expanded_key[752], expanded_key[753], expanded_key[754], expanded_key[755], expanded_key[756], expanded_key[757], expanded_key[758], expanded_key[759], expanded_key[760], expanded_key[761], expanded_key[762], expanded_key[763], expanded_key[764], expanded_key[765], expanded_key[766], expanded_key[767]};
        assign tmp1764 = mem_6[tmp1713];
    assign tmp1637 = tmp1635 ^ tmp1636;
    assign tmp1267 = {temp_19[8], temp_19[9], temp_19[10], temp_19[11], temp_19[12], temp_19[13], temp_19[14], temp_19[15]};
    assign tmp2343 = {temp_36[56], temp_36[57], temp_36[58], temp_36[59], temp_36[60], temp_36[61], temp_36[62], temp_36[63]};
    assign tmp137 = {tmp136[24], tmp136[25], tmp136[26], tmp136[27], tmp136[28], tmp136[29], tmp136[30], tmp136[31]};
        assign tmp1128 = mem_5[tmp1033];
    assign new_4 = tmp1712;
    assign tmp533 = tmp549;
        assign tmp1939 = mem_2[tmp1907];
        assign tmp326 = mem_2[tmp294];
    assign tmp617 = tmp615 ^ tmp616;
        assign tmp595 = mem_7[tmp563];
    assign tmp666 = {tmp665[0], tmp665[1], tmp665[2], tmp665[3], tmp665[4], tmp665[5], tmp665[6], tmp665[7]};
        assign tmp2026 = mem_6[tmp1947];
    assign tmp658 = {tmp657[0], tmp657[1], tmp657[2], tmp657[3], tmp657[4], tmp657[5], tmp657[6], tmp657[7]};
    assign tmp1974 = tmp2102;
    assign tmp420 = {tmp419[0], tmp419[1], tmp419[2], tmp419[3], tmp419[4], tmp419[5], tmp419[6], tmp419[7]};
    assign tmp1716 = {temp_27[96], temp_27[97], temp_27[98], temp_27[99], temp_27[100], temp_27[101], temp_27[102], temp_27[103]};
    assign tmp1339 = tmp1337 ^ tmp1338;
        assign tmp320 = mem_2[tmp288];
    assign shifted_w19 = tmp116;
    assign tmp305 = tmp321;
    assign tmp1030 = {temp_15[64], temp_15[65], temp_15[66], temp_15[67], temp_15[68], temp_15[69], temp_15[70], temp_15[71]};
    assign tmp1113 = tmp1111 ^ tmp1112;
    assign tmp15 = {tmp11[0], tmp11[1], tmp11[2], tmp11[3], tmp11[4], tmp11[5], tmp11[6], tmp11[7]};
    assign tmp265 = {new_state[120], new_state[121], new_state[122], new_state[123], new_state[124], new_state[125], new_state[126], new_state[127]};
        assign tmp1124 = mem_4[tmp1034];
    assign tmp2197 = tmp2276;
    assign tmp2284 = {tmp2283[0], tmp2283[1], tmp2283[2], tmp2283[3], tmp2283[4], tmp2283[5], tmp2283[6], tmp2283[7]};
    assign tmp671 = tmp669 ^ tmp670;
    assign tmp2009 = tmp2007 ^ tmp2008;
    assign b3_w39 = tmp244;
        assign tmp227 = mem_3[const226_9];
    assign tmp541 = tmp557;
    assign substituted_w19 = tmp125;
        assign tmp826 = mem_5[tmp794];
    assign tmp294 = {temp_1[24], temp_1[25], temp_1[26], temp_1[27], temp_1[28], temp_1[29], temp_1[30], temp_1[31]};
    assign tmp970 = {temp_12[0], temp_12[1], temp_12[2], temp_12[3], temp_12[4], temp_12[5], temp_12[6], temp_12[7]};
        assign tmp1143 = mem_7[tmp1034];
        assign tmp437 = mem_7[tmp342];
    assign tmp920 = {tmp919[0], tmp919[1], tmp919[2], tmp919[3], tmp919[4], tmp919[5], tmp919[6], tmp919[7]};
        assign tmp833 = mem_7[tmp794];
        assign tmp1614 = mem_6[tmp1497];
    assign tmp32 = concat_w3 ^ substituted_w3;
    assign tmp2054 = {tmp2053[0], tmp2053[1], tmp2053[2], tmp2053[3], tmp2053[4], tmp2053[5], tmp2053[6], tmp2053[7]};
        assign tmp1756 = mem_6[tmp1716];
        assign tmp1806 = mem_4[tmp1719];
    assign a4_w31 = tmp190;
        assign tmp667 = mem_7[tmp572];
    assign tmp1789 = tmp1787 ^ tmp1788;
        assign tmp2391 = mem_2[tmp2359];
        assign tmp402 = mem_4[tmp340];

    always @( posedge clk )
    begin
    end
endmodule


--- Verilog for the TestBench ---
module tb();
    reg clk;
    reg [127:0] aes_ciphertext;
    reg [127:0] aes_key;
    wire [127:0] aes_plaintext;

    toplevel block(.aes_plaintext(aes_plaintext), .aes_key(aes_key), .aes_ciphertext(aes_ciphertext), .clk(clk));

    always
        #0.5 clk = ~clk;

    initial begin
        $dumpfile ("waveform.vcd");
        $dumpvars;

        clk = 0;
        aes_ciphertext = 128'd136792598789324718765670228683992083246;
        aes_key = 128'd0;

        #2
        $finish;
    end
endmodule
